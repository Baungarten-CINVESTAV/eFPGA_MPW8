magic
tech sky130A
magscale 1 2
timestamp 1672417903
<< viali >>
rect 1593 37281 1627 37315
rect 9505 37281 9539 37315
rect 11713 37281 11747 37315
rect 22017 37281 22051 37315
rect 30941 37281 30975 37315
rect 34897 37281 34931 37315
rect 37473 37281 37507 37315
rect 1869 37213 1903 37247
rect 2881 37213 2915 37247
rect 4169 37213 4203 37247
rect 4813 37213 4847 37247
rect 6009 37213 6043 37247
rect 6745 37213 6779 37247
rect 7849 37213 7883 37247
rect 9781 37213 9815 37247
rect 11989 37213 12023 37247
rect 13185 37213 13219 37247
rect 14289 37213 14323 37247
rect 15761 37213 15795 37247
rect 17509 37213 17543 37247
rect 19625 37213 19659 37247
rect 20085 37213 20119 37247
rect 22293 37213 22327 37247
rect 24593 37213 24627 37247
rect 25513 37213 25547 37247
rect 27353 37213 27387 37247
rect 27813 37213 27847 37247
rect 28733 37213 28767 37247
rect 29929 37213 29963 37247
rect 31217 37213 31251 37247
rect 32321 37213 32355 37247
rect 33241 37213 33275 37247
rect 35173 37213 35207 37247
rect 36185 37213 36219 37247
rect 37749 37213 37783 37247
rect 3065 37077 3099 37111
rect 3985 37077 4019 37111
rect 4629 37077 4663 37111
rect 5825 37077 5859 37111
rect 6561 37077 6595 37111
rect 8033 37077 8067 37111
rect 9965 37077 9999 37111
rect 13001 37077 13035 37111
rect 14473 37077 14507 37111
rect 15577 37077 15611 37111
rect 17693 37077 17727 37111
rect 19441 37077 19475 37111
rect 20269 37077 20303 37111
rect 24777 37077 24811 37111
rect 25329 37077 25363 37111
rect 27169 37077 27203 37111
rect 27997 37077 28031 37111
rect 28549 37077 28583 37111
rect 29745 37077 29779 37111
rect 32505 37077 32539 37111
rect 33057 37077 33091 37111
rect 36369 37077 36403 37111
rect 9321 36873 9355 36907
rect 13185 36873 13219 36907
rect 17049 36873 17083 36907
rect 22201 36873 22235 36907
rect 26065 36873 26099 36907
rect 36829 36873 36863 36907
rect 38117 36805 38151 36839
rect 1593 36737 1627 36771
rect 3065 36737 3099 36771
rect 8861 36737 8895 36771
rect 9137 36737 9171 36771
rect 13369 36737 13403 36771
rect 14473 36737 14507 36771
rect 16865 36737 16899 36771
rect 22017 36737 22051 36771
rect 23305 36737 23339 36771
rect 26249 36737 26283 36771
rect 35541 36737 35575 36771
rect 36185 36737 36219 36771
rect 36645 36737 36679 36771
rect 1869 36669 1903 36703
rect 23581 36669 23615 36703
rect 14289 36601 14323 36635
rect 36001 36601 36035 36635
rect 2881 36533 2915 36567
rect 35357 36533 35391 36567
rect 38209 36533 38243 36567
rect 1777 36329 1811 36363
rect 35633 36329 35667 36363
rect 37473 36329 37507 36363
rect 36645 36261 36679 36295
rect 1593 36125 1627 36159
rect 2513 36125 2547 36159
rect 35541 36125 35575 36159
rect 36829 36125 36863 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 2329 35989 2363 36023
rect 38209 35989 38243 36023
rect 1593 35649 1627 35683
rect 38025 35649 38059 35683
rect 1777 35445 1811 35479
rect 38209 35445 38243 35479
rect 1777 35037 1811 35071
rect 37657 35037 37691 35071
rect 1593 34901 1627 34935
rect 37473 34901 37507 34935
rect 14197 34697 14231 34731
rect 35265 34697 35299 34731
rect 36001 34697 36035 34731
rect 14381 34561 14415 34595
rect 35449 34561 35483 34595
rect 35909 34561 35943 34595
rect 38025 34561 38059 34595
rect 38209 34357 38243 34391
rect 18981 33609 19015 33643
rect 1593 33473 1627 33507
rect 19165 33473 19199 33507
rect 1777 33337 1811 33371
rect 5733 32861 5767 32895
rect 23765 32861 23799 32895
rect 38025 32861 38059 32895
rect 5825 32725 5859 32759
rect 23857 32725 23891 32759
rect 38209 32725 38243 32759
rect 9045 32385 9079 32419
rect 38025 32385 38059 32419
rect 1593 32317 1627 32351
rect 1869 32317 1903 32351
rect 9137 32181 9171 32215
rect 38209 32181 38243 32215
rect 4537 31977 4571 32011
rect 7481 31977 7515 32011
rect 24685 31977 24719 32011
rect 9229 31909 9263 31943
rect 21833 31909 21867 31943
rect 15945 31841 15979 31875
rect 1593 31773 1627 31807
rect 4721 31773 4755 31807
rect 7665 31773 7699 31807
rect 9137 31773 9171 31807
rect 15853 31773 15887 31807
rect 21741 31773 21775 31807
rect 24593 31773 24627 31807
rect 1777 31637 1811 31671
rect 7481 31433 7515 31467
rect 7389 31297 7423 31331
rect 23949 31297 23983 31331
rect 28641 31297 28675 31331
rect 24041 31093 24075 31127
rect 28733 31093 28767 31127
rect 4997 30685 5031 30719
rect 9413 30685 9447 30719
rect 22109 30685 22143 30719
rect 38301 30685 38335 30719
rect 20085 30617 20119 30651
rect 20269 30617 20303 30651
rect 5089 30549 5123 30583
rect 9505 30549 9539 30583
rect 22201 30549 22235 30583
rect 38117 30549 38151 30583
rect 1593 30209 1627 30243
rect 12357 30209 12391 30243
rect 25881 30209 25915 30243
rect 27169 30209 27203 30243
rect 27261 30073 27295 30107
rect 1777 30005 1811 30039
rect 12449 30005 12483 30039
rect 25973 30005 26007 30039
rect 6745 29801 6779 29835
rect 6653 29597 6687 29631
rect 9137 29597 9171 29631
rect 38117 29529 38151 29563
rect 9229 29461 9263 29495
rect 38209 29461 38243 29495
rect 4445 29257 4479 29291
rect 33241 29257 33275 29291
rect 1777 29121 1811 29155
rect 4629 29121 4663 29155
rect 7113 29121 7147 29155
rect 33425 29121 33459 29155
rect 1593 28985 1627 29019
rect 7205 28985 7239 29019
rect 15117 28509 15151 28543
rect 26249 28509 26283 28543
rect 15209 28373 15243 28407
rect 26341 28373 26375 28407
rect 32321 28169 32355 28203
rect 17049 28101 17083 28135
rect 1777 28033 1811 28067
rect 18429 28033 18463 28067
rect 29285 28033 29319 28067
rect 29377 28033 29411 28067
rect 32505 28033 32539 28067
rect 38301 28033 38335 28067
rect 16957 27965 16991 27999
rect 17509 27897 17543 27931
rect 1593 27829 1627 27863
rect 18521 27829 18555 27863
rect 38117 27829 38151 27863
rect 28457 27557 28491 27591
rect 1593 27421 1627 27455
rect 2329 27421 2363 27455
rect 11621 27421 11655 27455
rect 12449 27421 12483 27455
rect 12909 27421 12943 27455
rect 13553 27421 13587 27455
rect 14289 27421 14323 27455
rect 28365 27421 28399 27455
rect 38025 27421 38059 27455
rect 1777 27285 1811 27319
rect 2421 27285 2455 27319
rect 11437 27285 11471 27319
rect 12265 27285 12299 27319
rect 13001 27285 13035 27319
rect 13645 27285 13679 27319
rect 14381 27285 14415 27319
rect 38209 27285 38243 27319
rect 5917 27081 5951 27115
rect 14565 27081 14599 27115
rect 6837 27013 6871 27047
rect 8769 27013 8803 27047
rect 9321 27013 9355 27047
rect 13461 27013 13495 27047
rect 1869 26945 1903 26979
rect 2513 26945 2547 26979
rect 3157 26945 3191 26979
rect 5825 26945 5859 26979
rect 6745 26945 6779 26979
rect 7941 26945 7975 26979
rect 11069 26945 11103 26979
rect 11713 26945 11747 26979
rect 12357 26945 12391 26979
rect 14473 26945 14507 26979
rect 32321 26945 32355 26979
rect 8677 26877 8711 26911
rect 13369 26877 13403 26911
rect 11805 26809 11839 26843
rect 13921 26809 13955 26843
rect 1961 26741 1995 26775
rect 2605 26741 2639 26775
rect 3249 26741 3283 26775
rect 8033 26741 8067 26775
rect 10885 26741 10919 26775
rect 12449 26741 12483 26775
rect 32413 26741 32447 26775
rect 18061 26537 18095 26571
rect 3985 26469 4019 26503
rect 6285 26469 6319 26503
rect 6929 26469 6963 26503
rect 10241 26469 10275 26503
rect 11345 26469 11379 26503
rect 38117 26469 38151 26503
rect 9873 26401 9907 26435
rect 10057 26401 10091 26435
rect 10977 26401 11011 26435
rect 14381 26401 14415 26435
rect 15393 26401 15427 26435
rect 16037 26401 16071 26435
rect 2053 26333 2087 26367
rect 2697 26333 2731 26367
rect 4169 26333 4203 26367
rect 6469 26333 6503 26367
rect 7113 26333 7147 26367
rect 11161 26333 11195 26367
rect 12265 26333 12299 26367
rect 18245 26333 18279 26367
rect 19625 26333 19659 26367
rect 20821 26333 20855 26367
rect 22385 26333 22419 26367
rect 23029 26333 23063 26367
rect 38301 26333 38335 26367
rect 2145 26265 2179 26299
rect 2789 26265 2823 26299
rect 14473 26265 14507 26299
rect 16129 26265 16163 26299
rect 17049 26265 17083 26299
rect 20913 26265 20947 26299
rect 12081 26197 12115 26231
rect 19441 26197 19475 26231
rect 22201 26197 22235 26231
rect 22845 26197 22879 26231
rect 16957 25993 16991 26027
rect 9505 25925 9539 25959
rect 18705 25925 18739 25959
rect 2145 25857 2179 25891
rect 3433 25857 3467 25891
rect 4077 25857 4111 25891
rect 4905 25857 4939 25891
rect 8033 25857 8067 25891
rect 9413 25857 9447 25891
rect 10793 25857 10827 25891
rect 12457 25855 12491 25889
rect 14105 25857 14139 25891
rect 16865 25857 16899 25891
rect 17969 25857 18003 25891
rect 19533 25857 19567 25891
rect 2789 25789 2823 25823
rect 7849 25789 7883 25823
rect 18061 25721 18095 25755
rect 2237 25653 2271 25687
rect 3525 25653 3559 25687
rect 4169 25653 4203 25687
rect 4721 25653 4755 25687
rect 8309 25653 8343 25687
rect 10885 25653 10919 25687
rect 12541 25653 12575 25687
rect 14197 25653 14231 25687
rect 18797 25653 18831 25687
rect 19349 25653 19383 25687
rect 5273 25449 5307 25483
rect 12817 25449 12851 25483
rect 32229 25449 32263 25483
rect 19717 25381 19751 25415
rect 1869 25313 1903 25347
rect 11345 25313 11379 25347
rect 12633 25313 12667 25347
rect 17141 25313 17175 25347
rect 17509 25313 17543 25347
rect 21557 25313 21591 25347
rect 1593 25245 1627 25279
rect 2881 25245 2915 25279
rect 3985 25245 4019 25279
rect 4629 25245 4663 25279
rect 5457 25245 5491 25279
rect 9597 25245 9631 25279
rect 10425 25245 10459 25279
rect 12449 25245 12483 25279
rect 18245 25245 18279 25279
rect 19533 25245 19567 25279
rect 20729 25245 20763 25279
rect 21373 25245 21407 25279
rect 27261 25245 27295 25279
rect 27353 25245 27387 25279
rect 32413 25245 32447 25279
rect 4077 25177 4111 25211
rect 11437 25177 11471 25211
rect 11989 25177 12023 25211
rect 17233 25177 17267 25211
rect 2973 25109 3007 25143
rect 4721 25109 4755 25143
rect 6837 25109 6871 25143
rect 9689 25109 9723 25143
rect 10517 25109 10551 25143
rect 16405 25109 16439 25143
rect 18337 25109 18371 25143
rect 22017 25109 22051 25143
rect 23581 24905 23615 24939
rect 6745 24837 6779 24871
rect 6837 24837 6871 24871
rect 8125 24837 8159 24871
rect 9321 24837 9355 24871
rect 14105 24837 14139 24871
rect 17049 24837 17083 24871
rect 17601 24837 17635 24871
rect 22201 24837 22235 24871
rect 2237 24769 2271 24803
rect 2697 24769 2731 24803
rect 3801 24769 3835 24803
rect 4629 24769 4663 24803
rect 5089 24769 5123 24803
rect 5917 24769 5951 24803
rect 11805 24769 11839 24803
rect 13277 24769 13311 24803
rect 15117 24769 15151 24803
rect 16129 24769 16163 24803
rect 16221 24769 16255 24803
rect 18061 24769 18095 24803
rect 18245 24769 18279 24803
rect 20177 24769 20211 24803
rect 23765 24769 23799 24803
rect 24409 24769 24443 24803
rect 29009 24769 29043 24803
rect 38025 24769 38059 24803
rect 8033 24701 8067 24735
rect 8309 24701 8343 24735
rect 9229 24701 9263 24735
rect 14013 24701 14047 24735
rect 16957 24701 16991 24735
rect 19993 24701 20027 24735
rect 20637 24701 20671 24735
rect 22109 24701 22143 24735
rect 5733 24633 5767 24667
rect 7297 24633 7331 24667
rect 9781 24633 9815 24667
rect 14565 24633 14599 24667
rect 22661 24633 22695 24667
rect 2053 24565 2087 24599
rect 2789 24565 2823 24599
rect 3893 24565 3927 24599
rect 4445 24565 4479 24599
rect 5181 24565 5215 24599
rect 11897 24565 11931 24599
rect 13369 24565 13403 24599
rect 15209 24565 15243 24599
rect 18705 24565 18739 24599
rect 24225 24565 24259 24599
rect 29101 24565 29135 24599
rect 38209 24565 38243 24599
rect 6193 24361 6227 24395
rect 23581 24361 23615 24395
rect 20913 24293 20947 24327
rect 8033 24225 8067 24259
rect 12541 24225 12575 24259
rect 13185 24225 13219 24259
rect 20361 24225 20395 24259
rect 1869 24157 1903 24191
rect 2513 24157 2547 24191
rect 4169 24157 4203 24191
rect 4997 24157 5031 24191
rect 5457 24157 5491 24191
rect 6101 24157 6135 24191
rect 7021 24157 7055 24191
rect 11161 24157 11195 24191
rect 14289 24157 14323 24191
rect 14933 24157 14967 24191
rect 16865 24157 16899 24191
rect 18153 24157 18187 24191
rect 19441 24157 19475 24191
rect 22845 24157 22879 24191
rect 23765 24157 23799 24191
rect 38025 24157 38059 24191
rect 2605 24089 2639 24123
rect 10057 24089 10091 24123
rect 10149 24089 10183 24123
rect 10701 24089 10735 24123
rect 12633 24089 12667 24123
rect 18245 24089 18279 24123
rect 20453 24089 20487 24123
rect 1961 24021 1995 24055
rect 3157 24021 3191 24055
rect 4261 24021 4295 24055
rect 4813 24021 4847 24055
rect 5549 24021 5583 24055
rect 7113 24021 7147 24055
rect 11253 24021 11287 24055
rect 14381 24021 14415 24055
rect 15025 24021 15059 24055
rect 16957 24021 16991 24055
rect 19533 24021 19567 24055
rect 22937 24021 22971 24055
rect 38209 24021 38243 24055
rect 7205 23817 7239 23851
rect 10977 23817 11011 23851
rect 19717 23817 19751 23851
rect 3341 23749 3375 23783
rect 8585 23749 8619 23783
rect 8677 23749 8711 23783
rect 12633 23749 12667 23783
rect 13737 23749 13771 23783
rect 13829 23749 13863 23783
rect 16037 23749 16071 23783
rect 17601 23749 17635 23783
rect 1869 23681 1903 23715
rect 4353 23681 4387 23715
rect 4997 23681 5031 23715
rect 5641 23681 5675 23715
rect 6561 23681 6595 23715
rect 7389 23681 7423 23715
rect 7849 23681 7883 23715
rect 9689 23681 9723 23715
rect 10517 23681 10551 23715
rect 11161 23681 11195 23715
rect 11805 23681 11839 23715
rect 14841 23681 14875 23715
rect 15945 23681 15979 23715
rect 19257 23681 19291 23715
rect 22569 23681 22603 23715
rect 23489 23681 23523 23715
rect 31217 23681 31251 23715
rect 2145 23613 2179 23647
rect 3249 23613 3283 23647
rect 7941 23613 7975 23647
rect 12541 23613 12575 23647
rect 13185 23613 13219 23647
rect 14933 23613 14967 23647
rect 17509 23613 17543 23647
rect 17969 23613 18003 23647
rect 19073 23613 19107 23647
rect 3801 23545 3835 23579
rect 6653 23545 6687 23579
rect 9137 23545 9171 23579
rect 14289 23545 14323 23579
rect 4445 23477 4479 23511
rect 5089 23477 5123 23511
rect 5733 23477 5767 23511
rect 9781 23477 9815 23511
rect 10333 23477 10367 23511
rect 11897 23477 11931 23511
rect 22661 23477 22695 23511
rect 23305 23477 23339 23511
rect 31309 23477 31343 23511
rect 3341 23273 3375 23307
rect 18337 23273 18371 23307
rect 30481 23273 30515 23307
rect 10517 23205 10551 23239
rect 4169 23137 4203 23171
rect 11161 23137 11195 23171
rect 11437 23137 11471 23171
rect 13093 23137 13127 23171
rect 16313 23137 16347 23171
rect 19533 23137 19567 23171
rect 3249 23069 3283 23103
rect 4077 23069 4111 23103
rect 4813 23069 4847 23103
rect 5825 23069 5859 23103
rect 6469 23069 6503 23103
rect 7113 23069 7147 23103
rect 7941 23069 7975 23103
rect 9229 23069 9263 23103
rect 12541 23069 12575 23103
rect 18521 23069 18555 23103
rect 23305 23069 23339 23103
rect 30665 23069 30699 23103
rect 1777 23001 1811 23035
rect 1869 23001 1903 23035
rect 2421 23001 2455 23035
rect 6561 23001 6595 23035
rect 9965 23001 9999 23035
rect 10057 23001 10091 23035
rect 11253 23001 11287 23035
rect 13185 23001 13219 23035
rect 13737 23001 13771 23035
rect 15117 23001 15151 23035
rect 15209 23001 15243 23035
rect 15761 23001 15795 23035
rect 16405 23001 16439 23035
rect 17325 23001 17359 23035
rect 19625 23001 19659 23035
rect 20177 23001 20211 23035
rect 4905 22933 4939 22967
rect 5917 22933 5951 22967
rect 7205 22933 7239 22967
rect 8033 22933 8067 22967
rect 9321 22933 9355 22967
rect 12357 22933 12391 22967
rect 14289 22933 14323 22967
rect 23121 22933 23155 22967
rect 4261 22729 4295 22763
rect 11805 22729 11839 22763
rect 1961 22661 1995 22695
rect 3065 22661 3099 22695
rect 3157 22661 3191 22695
rect 5181 22661 5215 22695
rect 10149 22661 10183 22695
rect 10701 22661 10735 22695
rect 12633 22661 12667 22695
rect 13185 22661 13219 22695
rect 13737 22661 13771 22695
rect 13829 22661 13863 22695
rect 16129 22661 16163 22695
rect 4169 22593 4203 22627
rect 5089 22593 5123 22627
rect 5825 22593 5859 22627
rect 5917 22593 5951 22627
rect 6837 22593 6871 22627
rect 7481 22593 7515 22627
rect 8677 22593 8711 22627
rect 9321 22593 9355 22627
rect 11713 22593 11747 22627
rect 15393 22593 15427 22627
rect 16037 22593 16071 22627
rect 18153 22593 18187 22627
rect 36737 22593 36771 22627
rect 38025 22593 38059 22627
rect 1869 22525 1903 22559
rect 2145 22525 2179 22559
rect 10057 22525 10091 22559
rect 12541 22525 12575 22559
rect 14381 22525 14415 22559
rect 3617 22457 3651 22491
rect 38209 22457 38243 22491
rect 2881 22389 2915 22423
rect 6929 22389 6963 22423
rect 7573 22389 7607 22423
rect 8769 22389 8803 22423
rect 9413 22389 9447 22423
rect 15485 22389 15519 22423
rect 18245 22389 18279 22423
rect 36829 22389 36863 22423
rect 37841 22185 37875 22219
rect 8493 22117 8527 22151
rect 18797 22117 18831 22151
rect 20637 22117 20671 22151
rect 6285 22049 6319 22083
rect 10241 22049 10275 22083
rect 15117 22049 15151 22083
rect 15945 22049 15979 22083
rect 17049 22049 17083 22083
rect 17325 22049 17359 22083
rect 18245 22049 18279 22083
rect 20085 22049 20119 22083
rect 25329 22049 25363 22083
rect 1593 21981 1627 22015
rect 1869 21981 1903 22015
rect 4261 21981 4295 22015
rect 4905 21981 4939 22015
rect 5549 21981 5583 22015
rect 6193 21981 6227 22015
rect 7113 21981 7147 22015
rect 7757 21981 7791 22015
rect 8425 21981 8459 22015
rect 12449 21981 12483 22015
rect 12909 21981 12943 22015
rect 13561 21975 13595 22009
rect 14381 21981 14415 22015
rect 38025 21981 38059 22015
rect 2973 21913 3007 21947
rect 4353 21913 4387 21947
rect 7205 21913 7239 21947
rect 9229 21913 9263 21947
rect 9321 21913 9355 21947
rect 10793 21913 10827 21947
rect 10885 21913 10919 21947
rect 11437 21913 11471 21947
rect 13645 21913 13679 21947
rect 15209 21913 15243 21947
rect 17141 21913 17175 21947
rect 18337 21913 18371 21947
rect 20177 21913 20211 21947
rect 25421 21913 25455 21947
rect 26341 21913 26375 21947
rect 3065 21845 3099 21879
rect 4997 21845 5031 21879
rect 5641 21845 5675 21879
rect 7849 21845 7883 21879
rect 12265 21845 12299 21879
rect 13001 21845 13035 21879
rect 14473 21845 14507 21879
rect 21741 21845 21775 21879
rect 5917 21641 5951 21675
rect 25237 21641 25271 21675
rect 32321 21641 32355 21675
rect 1869 21573 1903 21607
rect 3433 21573 3467 21607
rect 4629 21573 4663 21607
rect 7205 21573 7239 21607
rect 7297 21573 7331 21607
rect 8861 21573 8895 21607
rect 12173 21573 12207 21607
rect 13369 21573 13403 21607
rect 18521 21573 18555 21607
rect 19165 21573 19199 21607
rect 19901 21573 19935 21607
rect 25973 21573 26007 21607
rect 26065 21573 26099 21607
rect 5825 21505 5859 21539
rect 10333 21505 10367 21539
rect 10977 21505 11011 21539
rect 14381 21505 14415 21539
rect 15945 21505 15979 21539
rect 18429 21505 18463 21539
rect 19073 21505 19107 21539
rect 22017 21505 22051 21539
rect 22201 21505 22235 21539
rect 23765 21505 23799 21539
rect 25145 21505 25179 21539
rect 32505 21505 32539 21539
rect 38025 21505 38059 21539
rect 1777 21437 1811 21471
rect 2789 21437 2823 21471
rect 3341 21437 3375 21471
rect 3801 21437 3835 21471
rect 4537 21437 4571 21471
rect 7481 21437 7515 21471
rect 8769 21437 8803 21471
rect 9045 21437 9079 21471
rect 12081 21437 12115 21471
rect 13277 21437 13311 21471
rect 14565 21437 14599 21471
rect 19809 21437 19843 21471
rect 23121 21437 23155 21471
rect 23305 21437 23339 21471
rect 5089 21369 5123 21403
rect 12633 21369 12667 21403
rect 13829 21369 13863 21403
rect 15025 21369 15059 21403
rect 20361 21369 20395 21403
rect 26525 21369 26559 21403
rect 10425 21301 10459 21335
rect 11069 21301 11103 21335
rect 16037 21301 16071 21335
rect 22385 21301 22419 21335
rect 38209 21301 38243 21335
rect 9413 21097 9447 21131
rect 16129 21097 16163 21131
rect 20545 21097 20579 21131
rect 26249 21097 26283 21131
rect 29837 21097 29871 21131
rect 32597 21097 32631 21131
rect 5273 21029 5307 21063
rect 23949 21029 23983 21063
rect 2237 20961 2271 20995
rect 2881 20961 2915 20995
rect 6561 20961 6595 20995
rect 10057 20961 10091 20995
rect 10977 20961 11011 20995
rect 12541 20961 12575 20995
rect 14657 20961 14691 20995
rect 17233 20961 17267 20995
rect 17509 20961 17543 20995
rect 3985 20893 4019 20927
rect 9321 20893 9355 20927
rect 11805 20893 11839 20927
rect 15669 20893 15703 20927
rect 16313 20893 16347 20927
rect 20453 20893 20487 20927
rect 25513 20893 25547 20927
rect 26157 20893 26191 20927
rect 26985 20893 27019 20927
rect 29745 20893 29779 20927
rect 32781 20893 32815 20927
rect 37473 20893 37507 20927
rect 37749 20893 37783 20927
rect 2329 20825 2363 20859
rect 4721 20825 4755 20859
rect 4813 20825 4847 20859
rect 5917 20825 5951 20859
rect 6009 20825 6043 20859
rect 7481 20825 7515 20859
rect 7573 20825 7607 20859
rect 8125 20825 8159 20859
rect 10149 20825 10183 20859
rect 12633 20825 12667 20859
rect 13553 20825 13587 20859
rect 14381 20825 14415 20859
rect 14473 20825 14507 20859
rect 17325 20825 17359 20859
rect 23397 20825 23431 20859
rect 23489 20825 23523 20859
rect 25605 20825 25639 20859
rect 4077 20757 4111 20791
rect 11897 20757 11931 20791
rect 15485 20757 15519 20791
rect 24869 20757 24903 20791
rect 26801 20757 26835 20791
rect 17601 20553 17635 20587
rect 23673 20553 23707 20587
rect 24225 20553 24259 20587
rect 1685 20485 1719 20519
rect 1777 20485 1811 20519
rect 2697 20485 2731 20519
rect 3341 20485 3375 20519
rect 3893 20485 3927 20519
rect 4537 20485 4571 20519
rect 5089 20485 5123 20519
rect 6653 20485 6687 20519
rect 6745 20485 6779 20519
rect 8217 20485 8251 20519
rect 10517 20485 10551 20519
rect 10609 20485 10643 20519
rect 11897 20485 11931 20519
rect 12817 20485 12851 20519
rect 13818 20485 13852 20519
rect 13930 20485 13964 20519
rect 14841 20485 14875 20519
rect 15485 20485 15519 20519
rect 18521 20485 18555 20519
rect 25789 20485 25823 20519
rect 5825 20417 5859 20451
rect 16957 20417 16991 20451
rect 17141 20417 17175 20451
rect 23581 20417 23615 20451
rect 24409 20417 24443 20451
rect 3249 20349 3283 20383
rect 4445 20349 4479 20383
rect 6929 20349 6963 20383
rect 8125 20349 8159 20383
rect 9137 20349 9171 20383
rect 9781 20349 9815 20383
rect 11805 20349 11839 20383
rect 15393 20349 15427 20383
rect 15669 20349 15703 20383
rect 18429 20349 18463 20383
rect 19441 20349 19475 20383
rect 25697 20349 25731 20383
rect 26341 20349 26375 20383
rect 11069 20281 11103 20315
rect 5917 20213 5951 20247
rect 16405 20009 16439 20043
rect 18153 20009 18187 20043
rect 25789 20009 25823 20043
rect 2421 19873 2455 19907
rect 3433 19873 3467 19907
rect 5089 19873 5123 19907
rect 7849 19873 7883 19907
rect 9597 19873 9631 19907
rect 10517 19873 10551 19907
rect 12081 19873 12115 19907
rect 13553 19873 13587 19907
rect 14381 19873 14415 19907
rect 21741 19873 21775 19907
rect 23397 19873 23431 19907
rect 24041 19873 24075 19907
rect 1777 19805 1811 19839
rect 4353 19805 4387 19839
rect 6837 19805 6871 19839
rect 16313 19805 16347 19839
rect 17049 19805 17083 19839
rect 18061 19805 18095 19839
rect 22569 19805 22603 19839
rect 24593 19805 24627 19839
rect 25973 19805 26007 19839
rect 32045 19805 32079 19839
rect 2513 19737 2547 19771
rect 5181 19737 5215 19771
rect 6101 19737 6135 19771
rect 7021 19737 7055 19771
rect 7573 19737 7607 19771
rect 7665 19737 7699 19771
rect 9321 19737 9355 19771
rect 9413 19737 9447 19771
rect 10609 19737 10643 19771
rect 11529 19737 11563 19771
rect 12173 19737 12207 19771
rect 13093 19737 13127 19771
rect 14473 19737 14507 19771
rect 15393 19737 15427 19771
rect 21465 19737 21499 19771
rect 21557 19737 21591 19771
rect 23489 19737 23523 19771
rect 1777 19669 1811 19703
rect 4445 19669 4479 19703
rect 17141 19669 17175 19703
rect 22661 19669 22695 19703
rect 24685 19669 24719 19703
rect 32137 19669 32171 19703
rect 6837 19465 6871 19499
rect 16957 19465 16991 19499
rect 23949 19465 23983 19499
rect 30021 19465 30055 19499
rect 38117 19465 38151 19499
rect 1685 19397 1719 19431
rect 1777 19397 1811 19431
rect 2697 19397 2731 19431
rect 10241 19397 10275 19431
rect 12173 19397 12207 19431
rect 12909 19397 12943 19431
rect 14197 19397 14231 19431
rect 14289 19397 14323 19431
rect 15761 19397 15795 19431
rect 17969 19397 18003 19431
rect 18889 19397 18923 19431
rect 20085 19397 20119 19431
rect 24961 19397 24995 19431
rect 25513 19397 25547 19431
rect 3249 19329 3283 19363
rect 3985 19329 4019 19363
rect 6745 19329 6779 19363
rect 12081 19329 12115 19363
rect 15669 19329 15703 19363
rect 16865 19329 16899 19363
rect 21465 19329 21499 19363
rect 22201 19329 22235 19363
rect 23397 19329 23431 19363
rect 23857 19329 23891 19363
rect 29929 19329 29963 19363
rect 38301 19329 38335 19363
rect 5733 19261 5767 19295
rect 7389 19261 7423 19295
rect 7665 19261 7699 19295
rect 10149 19261 10183 19295
rect 11069 19261 11103 19295
rect 12817 19261 12851 19295
rect 13461 19261 13495 19295
rect 14657 19261 14691 19295
rect 17877 19261 17911 19295
rect 24869 19261 24903 19295
rect 25973 19261 26007 19295
rect 22017 19193 22051 19227
rect 3341 19125 3375 19159
rect 4248 19125 4282 19159
rect 9137 19125 9171 19159
rect 20177 19125 20211 19159
rect 21281 19125 21315 19159
rect 23213 19125 23247 19159
rect 3341 18921 3375 18955
rect 3985 18921 4019 18955
rect 8585 18921 8619 18955
rect 15577 18921 15611 18955
rect 17233 18921 17267 18955
rect 19717 18921 19751 18955
rect 25329 18921 25363 18955
rect 26065 18853 26099 18887
rect 1869 18785 1903 18819
rect 15025 18785 15059 18819
rect 23673 18785 23707 18819
rect 24961 18785 24995 18819
rect 25145 18785 25179 18819
rect 1593 18717 1627 18751
rect 4169 18717 4203 18751
rect 6837 18717 6871 18751
rect 9321 18717 9355 18751
rect 9965 18717 9999 18751
rect 12173 18717 12207 18751
rect 13277 18717 13311 18751
rect 15485 18717 15519 18751
rect 16497 18717 16531 18751
rect 17141 18717 17175 18751
rect 19625 18717 19659 18751
rect 20269 18717 20303 18751
rect 26249 18717 26283 18751
rect 4445 18649 4479 18683
rect 7113 18649 7147 18683
rect 10701 18649 10735 18683
rect 10793 18649 10827 18683
rect 11713 18649 11747 18683
rect 13553 18649 13587 18683
rect 14381 18649 14415 18683
rect 14473 18649 14507 18683
rect 23029 18649 23063 18683
rect 23121 18649 23155 18683
rect 5917 18581 5951 18615
rect 9413 18581 9447 18615
rect 10057 18581 10091 18615
rect 12265 18581 12299 18615
rect 16589 18581 16623 18615
rect 20361 18581 20395 18615
rect 3341 18377 3375 18411
rect 23213 18377 23247 18411
rect 23857 18377 23891 18411
rect 25053 18377 25087 18411
rect 8585 18309 8619 18343
rect 9321 18309 9355 18343
rect 11989 18309 12023 18343
rect 14197 18309 14231 18343
rect 19073 18309 19107 18343
rect 19165 18309 19199 18343
rect 4077 18241 4111 18275
rect 6561 18241 6595 18275
rect 9045 18241 9079 18275
rect 15761 18241 15795 18275
rect 18061 18241 18095 18275
rect 23397 18241 23431 18275
rect 24041 18241 24075 18275
rect 25237 18241 25271 18275
rect 25697 18241 25731 18275
rect 35357 18241 35391 18275
rect 38025 18241 38059 18275
rect 1593 18173 1627 18207
rect 1869 18173 1903 18207
rect 4353 18173 4387 18207
rect 5825 18173 5859 18207
rect 6837 18173 6871 18207
rect 11713 18173 11747 18207
rect 14105 18173 14139 18207
rect 15117 18173 15151 18207
rect 15577 18173 15611 18207
rect 19349 18173 19383 18207
rect 10793 18037 10827 18071
rect 13461 18037 13495 18071
rect 16221 18037 16255 18071
rect 18153 18037 18187 18071
rect 25789 18037 25823 18071
rect 35173 18037 35207 18071
rect 38209 18037 38243 18071
rect 15945 17833 15979 17867
rect 3433 17765 3467 17799
rect 1685 17697 1719 17731
rect 4077 17697 4111 17731
rect 6837 17697 6871 17731
rect 8585 17697 8619 17731
rect 9137 17697 9171 17731
rect 11621 17697 11655 17731
rect 13369 17697 13403 17731
rect 14381 17697 14415 17731
rect 19717 17697 19751 17731
rect 20821 17697 20855 17731
rect 21005 17697 21039 17731
rect 15853 17629 15887 17663
rect 16497 17629 16531 17663
rect 17141 17629 17175 17663
rect 1961 17561 1995 17595
rect 4353 17561 4387 17595
rect 7113 17561 7147 17595
rect 9413 17561 9447 17595
rect 11161 17561 11195 17595
rect 11897 17561 11931 17595
rect 14473 17561 14507 17595
rect 15393 17561 15427 17595
rect 19809 17561 19843 17595
rect 20361 17561 20395 17595
rect 5825 17493 5859 17527
rect 16589 17493 16623 17527
rect 17233 17493 17267 17527
rect 21465 17493 21499 17527
rect 6009 17289 6043 17323
rect 16957 17289 16991 17323
rect 34253 17289 34287 17323
rect 1869 17221 1903 17255
rect 4537 17221 4571 17255
rect 10793 17221 10827 17255
rect 11989 17221 12023 17255
rect 14197 17221 14231 17255
rect 15669 17221 15703 17255
rect 15761 17221 15795 17255
rect 23121 17221 23155 17255
rect 24501 17221 24535 17255
rect 6653 17153 6687 17187
rect 10057 17153 10091 17187
rect 11713 17153 11747 17187
rect 16865 17153 16899 17187
rect 17877 17153 17911 17187
rect 20085 17153 20119 17187
rect 23673 17153 23707 17187
rect 34437 17153 34471 17187
rect 1593 17085 1627 17119
rect 3617 17085 3651 17119
rect 4261 17085 4295 17119
rect 7757 17085 7791 17119
rect 8033 17085 8067 17119
rect 13737 17085 13771 17119
rect 14933 17085 14967 17119
rect 23029 17085 23063 17119
rect 24409 17085 24443 17119
rect 25421 17085 25455 17119
rect 16221 17017 16255 17051
rect 6745 16949 6779 16983
rect 9505 16949 9539 16983
rect 17969 16949 18003 16983
rect 20177 16949 20211 16983
rect 5720 16745 5754 16779
rect 9321 16745 9355 16779
rect 10609 16745 10643 16779
rect 11424 16745 11458 16779
rect 13645 16745 13679 16779
rect 16037 16745 16071 16779
rect 12909 16677 12943 16711
rect 1685 16609 1719 16643
rect 1961 16609 1995 16643
rect 5457 16609 5491 16643
rect 8401 16609 8435 16643
rect 11161 16609 11195 16643
rect 16681 16609 16715 16643
rect 18337 16609 18371 16643
rect 24685 16609 24719 16643
rect 26157 16609 26191 16643
rect 26341 16609 26375 16643
rect 9221 16551 9255 16585
rect 9873 16541 9907 16575
rect 9965 16541 9999 16575
rect 10517 16541 10551 16575
rect 13553 16541 13587 16575
rect 14749 16541 14783 16575
rect 15945 16541 15979 16575
rect 18153 16541 18187 16575
rect 19901 16541 19935 16575
rect 20821 16541 20855 16575
rect 23121 16541 23155 16575
rect 23857 16541 23891 16575
rect 23949 16541 23983 16575
rect 27813 16541 27847 16575
rect 27905 16541 27939 16575
rect 38025 16541 38059 16575
rect 3985 16473 4019 16507
rect 4721 16473 4755 16507
rect 7665 16473 7699 16507
rect 15025 16473 15059 16507
rect 16773 16473 16807 16507
rect 17693 16473 17727 16507
rect 18797 16473 18831 16507
rect 24777 16473 24811 16507
rect 25697 16473 25731 16507
rect 3433 16405 3467 16439
rect 7205 16405 7239 16439
rect 19993 16405 20027 16439
rect 20637 16405 20671 16439
rect 23213 16405 23247 16439
rect 26801 16405 26835 16439
rect 38209 16405 38243 16439
rect 3525 16201 3559 16235
rect 6009 16201 6043 16235
rect 10609 16201 10643 16235
rect 14381 16201 14415 16235
rect 20821 16201 20855 16235
rect 26341 16201 26375 16235
rect 27721 16201 27755 16235
rect 28273 16201 28307 16235
rect 7389 16133 7423 16167
rect 15761 16133 15795 16167
rect 17049 16133 17083 16167
rect 19441 16133 19475 16167
rect 22201 16133 22235 16167
rect 1777 16065 1811 16099
rect 4261 16065 4295 16099
rect 7113 16065 7147 16099
rect 9137 16065 9171 16099
rect 9873 16065 9907 16099
rect 10517 16065 10551 16099
rect 14289 16065 14323 16099
rect 14933 16065 14967 16099
rect 15669 16065 15703 16099
rect 21005 16065 21039 16099
rect 26249 16065 26283 16099
rect 27629 16065 27663 16099
rect 28457 16065 28491 16099
rect 29101 16065 29135 16099
rect 38025 16065 38059 16099
rect 2053 15997 2087 16031
rect 4537 15997 4571 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 15025 15997 15059 16031
rect 16957 15997 16991 16031
rect 18613 15997 18647 16031
rect 19349 15997 19383 16031
rect 20269 15997 20303 16031
rect 22109 15997 22143 16031
rect 22385 15997 22419 16031
rect 24225 15997 24259 16031
rect 9965 15929 9999 15963
rect 17509 15929 17543 15963
rect 13461 15861 13495 15895
rect 28917 15861 28951 15895
rect 38209 15861 38243 15895
rect 3341 15657 3375 15691
rect 4248 15657 4282 15691
rect 11805 15657 11839 15691
rect 22477 15657 22511 15691
rect 25237 15657 25271 15691
rect 5733 15589 5767 15623
rect 15577 15589 15611 15623
rect 22937 15589 22971 15623
rect 1593 15521 1627 15555
rect 1869 15521 1903 15555
rect 6561 15521 6595 15555
rect 10057 15521 10091 15555
rect 24593 15521 24627 15555
rect 24777 15521 24811 15555
rect 3985 15453 4019 15487
rect 9413 15453 9447 15487
rect 14841 15453 14875 15487
rect 15485 15453 15519 15487
rect 16129 15453 16163 15487
rect 17233 15453 17267 15487
rect 17325 15453 17359 15487
rect 17877 15453 17911 15487
rect 18521 15453 18555 15487
rect 21833 15453 21867 15487
rect 22017 15453 22051 15487
rect 23121 15453 23155 15487
rect 23765 15453 23799 15487
rect 28733 15453 28767 15487
rect 6837 15385 6871 15419
rect 10333 15385 10367 15419
rect 12725 15385 12759 15419
rect 12817 15385 12851 15419
rect 13737 15385 13771 15419
rect 19533 15385 19567 15419
rect 19625 15385 19659 15419
rect 20177 15385 20211 15419
rect 21189 15385 21223 15419
rect 8309 15317 8343 15351
rect 9505 15317 9539 15351
rect 14933 15317 14967 15351
rect 16221 15317 16255 15351
rect 17969 15317 18003 15351
rect 18613 15317 18647 15351
rect 21281 15317 21315 15351
rect 23581 15317 23615 15351
rect 28549 15317 28583 15351
rect 11069 15113 11103 15147
rect 13461 15113 13495 15147
rect 18521 15113 18555 15147
rect 20729 15113 20763 15147
rect 22109 15113 22143 15147
rect 1869 15045 1903 15079
rect 4261 15045 4295 15079
rect 10057 15045 10091 15079
rect 14197 15045 14231 15079
rect 15117 15045 15151 15079
rect 17049 15045 17083 15079
rect 19901 15045 19935 15079
rect 24133 15045 24167 15079
rect 1593 14977 1627 15011
rect 3985 14977 4019 15011
rect 6929 14977 6963 15011
rect 7389 14977 7423 15011
rect 10977 14977 11011 15011
rect 18429 14977 18463 15011
rect 19441 14977 19475 15011
rect 20637 14977 20671 15011
rect 21281 14977 21315 15011
rect 22017 14977 22051 15011
rect 24041 14977 24075 15011
rect 26249 14977 26283 15011
rect 28825 14977 28859 15011
rect 38025 14977 38059 15011
rect 3341 14909 3375 14943
rect 5733 14909 5767 14943
rect 8033 14909 8067 14943
rect 8309 14909 8343 14943
rect 11713 14909 11747 14943
rect 11989 14909 12023 14943
rect 14105 14909 14139 14943
rect 16129 14909 16163 14943
rect 16957 14909 16991 14943
rect 17601 14909 17635 14943
rect 19257 14909 19291 14943
rect 21373 14909 21407 14943
rect 27169 14909 27203 14943
rect 27353 14909 27387 14943
rect 6745 14841 6779 14875
rect 28641 14841 28675 14875
rect 7481 14773 7515 14807
rect 26341 14773 26375 14807
rect 27537 14773 27571 14807
rect 37841 14773 37875 14807
rect 4905 14569 4939 14603
rect 7205 14569 7239 14603
rect 7849 14569 7883 14603
rect 14657 14569 14691 14603
rect 20637 14569 20671 14603
rect 35357 14569 35391 14603
rect 13369 14501 13403 14535
rect 20085 14501 20119 14535
rect 1593 14433 1627 14467
rect 3341 14433 3375 14467
rect 4169 14433 4203 14467
rect 5733 14433 5767 14467
rect 9137 14433 9171 14467
rect 15485 14433 15519 14467
rect 15761 14433 15795 14467
rect 17417 14433 17451 14467
rect 19441 14433 19475 14467
rect 19625 14433 19659 14467
rect 24593 14433 24627 14467
rect 24777 14433 24811 14467
rect 26709 14433 26743 14467
rect 4813 14365 4847 14399
rect 5457 14365 5491 14399
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 11161 14365 11195 14399
rect 11621 14365 11655 14399
rect 14565 14365 14599 14399
rect 18705 14365 18739 14399
rect 20545 14365 20579 14399
rect 21741 14365 21775 14399
rect 27537 14365 27571 14399
rect 27997 14365 28031 14399
rect 35541 14365 35575 14399
rect 38025 14365 38059 14399
rect 1869 14297 1903 14331
rect 8493 14297 8527 14331
rect 9413 14297 9447 14331
rect 11897 14297 11931 14331
rect 15577 14297 15611 14331
rect 17509 14297 17543 14331
rect 18061 14297 18095 14331
rect 18797 14229 18831 14263
rect 21833 14229 21867 14263
rect 25237 14229 25271 14263
rect 27353 14229 27387 14263
rect 28089 14229 28123 14263
rect 38209 14229 38243 14263
rect 1777 14025 1811 14059
rect 13461 14025 13495 14059
rect 15669 14025 15703 14059
rect 26617 14025 26651 14059
rect 27169 14025 27203 14059
rect 33701 14025 33735 14059
rect 2421 13957 2455 13991
rect 6653 13957 6687 13991
rect 9873 13957 9907 13991
rect 10425 13957 10459 13991
rect 11069 13957 11103 13991
rect 14105 13957 14139 13991
rect 17049 13957 17083 13991
rect 17141 13957 17175 13991
rect 18061 13957 18095 13991
rect 18705 13957 18739 13991
rect 20361 13957 20395 13991
rect 1593 13889 1627 13923
rect 2237 13889 2271 13923
rect 2789 13889 2823 13923
rect 3065 13889 3099 13923
rect 6561 13889 6595 13923
rect 7205 13889 7239 13923
rect 10333 13889 10367 13923
rect 10977 13889 11011 13923
rect 11713 13889 11747 13923
rect 15577 13889 15611 13923
rect 20821 13889 20855 13923
rect 22937 13889 22971 13923
rect 23581 13889 23615 13923
rect 25973 13889 26007 13923
rect 26157 13889 26191 13923
rect 27353 13889 27387 13923
rect 27813 13889 27847 13923
rect 27905 13889 27939 13923
rect 33885 13889 33919 13923
rect 4261 13821 4295 13855
rect 4537 13821 4571 13855
rect 6009 13821 6043 13855
rect 7849 13821 7883 13855
rect 8125 13821 8159 13855
rect 11989 13821 12023 13855
rect 14013 13821 14047 13855
rect 15025 13821 15059 13855
rect 18613 13821 18647 13855
rect 18889 13821 18923 13855
rect 19717 13821 19751 13855
rect 19901 13821 19935 13855
rect 20913 13821 20947 13855
rect 22293 13821 22327 13855
rect 22477 13821 22511 13855
rect 3249 13685 3283 13719
rect 7297 13685 7331 13719
rect 23397 13685 23431 13719
rect 1856 13481 1890 13515
rect 3341 13481 3375 13515
rect 10885 13481 10919 13515
rect 19901 13481 19935 13515
rect 21649 13481 21683 13515
rect 22477 13481 22511 13515
rect 26801 13481 26835 13515
rect 7573 13413 7607 13447
rect 1593 13345 1627 13379
rect 9137 13345 9171 13379
rect 11345 13345 11379 13379
rect 14381 13345 14415 13379
rect 15393 13345 15427 13379
rect 16589 13345 16623 13379
rect 16957 13345 16991 13379
rect 20637 13345 20671 13379
rect 21097 13345 21131 13379
rect 3985 13277 4019 13311
rect 5825 13277 5859 13311
rect 8401 13277 8435 13311
rect 13369 13277 13403 13311
rect 15853 13277 15887 13311
rect 18613 13277 18647 13311
rect 19809 13277 19843 13311
rect 20453 13277 20487 13311
rect 21557 13277 21591 13311
rect 22661 13277 22695 13311
rect 23949 13277 23983 13311
rect 26157 13277 26191 13311
rect 26341 13277 26375 13311
rect 27261 13277 27295 13311
rect 38025 13277 38059 13311
rect 4721 13209 4755 13243
rect 6101 13209 6135 13243
rect 9413 13209 9447 13243
rect 11621 13209 11655 13243
rect 14473 13209 14507 13243
rect 16681 13209 16715 13243
rect 17877 13209 17911 13243
rect 8493 13141 8527 13175
rect 15945 13141 15979 13175
rect 17969 13141 18003 13175
rect 18705 13141 18739 13175
rect 23765 13141 23799 13175
rect 27353 13141 27387 13175
rect 38209 13141 38243 13175
rect 6009 12937 6043 12971
rect 6653 12937 6687 12971
rect 1869 12869 1903 12903
rect 9229 12869 9263 12903
rect 9689 12869 9723 12903
rect 13737 12869 13771 12903
rect 14197 12869 14231 12903
rect 15761 12869 15795 12903
rect 18705 12869 18739 12903
rect 22753 12869 22787 12903
rect 23397 12869 23431 12903
rect 6561 12801 6595 12835
rect 7205 12801 7239 12835
rect 11713 12801 11747 12835
rect 17233 12801 17267 12835
rect 17877 12801 17911 12835
rect 20085 12801 20119 12835
rect 20729 12801 20763 12835
rect 22017 12801 22051 12835
rect 22661 12801 22695 12835
rect 23305 12801 23339 12835
rect 38301 12801 38335 12835
rect 1593 12733 1627 12767
rect 3341 12733 3375 12767
rect 4261 12733 4295 12767
rect 4537 12733 4571 12767
rect 7481 12733 7515 12767
rect 10517 12733 10551 12767
rect 11989 12733 12023 12767
rect 14933 12733 14967 12767
rect 15669 12733 15703 12767
rect 18613 12733 18647 12767
rect 19625 12733 19659 12767
rect 16221 12665 16255 12699
rect 17325 12597 17359 12631
rect 17969 12597 18003 12631
rect 20177 12597 20211 12631
rect 20821 12597 20855 12631
rect 22109 12597 22143 12631
rect 38117 12597 38151 12631
rect 8493 12393 8527 12427
rect 13001 12393 13035 12427
rect 13553 12393 13587 12427
rect 22661 12393 22695 12427
rect 23305 12393 23339 12427
rect 16037 12325 16071 12359
rect 19901 12325 19935 12359
rect 1685 12257 1719 12291
rect 7021 12257 7055 12291
rect 9873 12257 9907 12291
rect 11253 12257 11287 12291
rect 17693 12257 17727 12291
rect 17877 12257 17911 12291
rect 22017 12257 22051 12291
rect 3985 12189 4019 12223
rect 6745 12189 6779 12223
rect 10609 12189 10643 12223
rect 13737 12189 13771 12223
rect 14289 12189 14323 12223
rect 18337 12189 18371 12223
rect 21925 12189 21959 12223
rect 22569 12189 22603 12223
rect 23213 12189 23247 12223
rect 23857 12189 23891 12223
rect 29745 12189 29779 12223
rect 1961 12121 1995 12155
rect 4261 12121 4295 12155
rect 9137 12121 9171 12155
rect 11529 12121 11563 12155
rect 14565 12121 14599 12155
rect 16589 12121 16623 12155
rect 16681 12121 16715 12155
rect 17233 12121 17267 12155
rect 19717 12121 19751 12155
rect 20453 12121 20487 12155
rect 20545 12121 20579 12155
rect 21465 12121 21499 12155
rect 29837 12121 29871 12155
rect 3433 12053 3467 12087
rect 5733 12053 5767 12087
rect 10701 12053 10735 12087
rect 23949 12053 23983 12087
rect 10425 11849 10459 11883
rect 15761 11849 15795 11883
rect 24869 11849 24903 11883
rect 1869 11781 1903 11815
rect 11989 11781 12023 11815
rect 14289 11781 14323 11815
rect 17049 11781 17083 11815
rect 19073 11781 19107 11815
rect 20545 11781 20579 11815
rect 22201 11781 22235 11815
rect 23121 11781 23155 11815
rect 1593 11713 1627 11747
rect 4261 11713 4295 11747
rect 6653 11713 6687 11747
rect 7297 11713 7331 11747
rect 7941 11713 7975 11747
rect 10333 11713 10367 11747
rect 10977 11713 11011 11747
rect 11713 11713 11747 11747
rect 14013 11713 14047 11747
rect 24133 11713 24167 11747
rect 24777 11713 24811 11747
rect 25697 11713 25731 11747
rect 29653 11713 29687 11747
rect 3617 11645 3651 11679
rect 4537 11645 4571 11679
rect 6745 11645 6779 11679
rect 8217 11645 8251 11679
rect 13461 11645 13495 11679
rect 16957 11645 16991 11679
rect 17233 11645 17267 11679
rect 18245 11645 18279 11679
rect 18981 11645 19015 11679
rect 20453 11645 20487 11679
rect 21373 11645 21407 11679
rect 22109 11645 22143 11679
rect 19533 11577 19567 11611
rect 6009 11509 6043 11543
rect 7389 11509 7423 11543
rect 9689 11509 9723 11543
rect 11069 11509 11103 11543
rect 24225 11509 24259 11543
rect 25513 11509 25547 11543
rect 29745 11509 29779 11543
rect 6101 11305 6135 11339
rect 6916 11305 6950 11339
rect 8401 11305 8435 11339
rect 9965 11305 9999 11339
rect 10609 11305 10643 11339
rect 38117 11305 38151 11339
rect 9321 11237 9355 11271
rect 12909 11237 12943 11271
rect 13645 11237 13679 11271
rect 1593 11169 1627 11203
rect 3341 11169 3375 11203
rect 4353 11169 4387 11203
rect 6653 11169 6687 11203
rect 16037 11169 16071 11203
rect 16589 11169 16623 11203
rect 18245 11169 18279 11203
rect 20177 11169 20211 11203
rect 9229 11101 9263 11135
rect 9873 11101 9907 11135
rect 10517 11101 10551 11135
rect 11161 11101 11195 11135
rect 13553 11101 13587 11135
rect 14289 11101 14323 11135
rect 18061 11101 18095 11135
rect 19441 11101 19475 11135
rect 23305 11101 23339 11135
rect 24777 11101 24811 11135
rect 26157 11101 26191 11135
rect 38301 11101 38335 11135
rect 1869 11033 1903 11067
rect 4629 11033 4663 11067
rect 11437 11033 11471 11067
rect 14565 11033 14599 11067
rect 16681 11033 16715 11067
rect 17601 11033 17635 11067
rect 19533 11033 19567 11067
rect 20269 11033 20303 11067
rect 21189 11033 21223 11067
rect 21833 11033 21867 11067
rect 21925 11033 21959 11067
rect 22845 11033 22879 11067
rect 23397 10965 23431 10999
rect 24593 10965 24627 10999
rect 25973 10965 26007 10999
rect 26617 10965 26651 10999
rect 1777 10761 1811 10795
rect 2329 10761 2363 10795
rect 3065 10761 3099 10795
rect 3709 10761 3743 10795
rect 6009 10761 6043 10795
rect 7297 10761 7331 10795
rect 11069 10761 11103 10795
rect 23581 10761 23615 10795
rect 24133 10761 24167 10795
rect 4537 10693 4571 10727
rect 8125 10693 8159 10727
rect 14289 10693 14323 10727
rect 18521 10693 18555 10727
rect 19441 10693 19475 10727
rect 20269 10693 20303 10727
rect 21189 10693 21223 10727
rect 29377 10693 29411 10727
rect 1685 10625 1719 10659
rect 2513 10625 2547 10659
rect 2973 10625 3007 10659
rect 3617 10625 3651 10659
rect 4261 10625 4295 10659
rect 6561 10625 6595 10659
rect 7205 10625 7239 10659
rect 7849 10625 7883 10659
rect 10333 10625 10367 10659
rect 10977 10625 11011 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 22385 10625 22419 10659
rect 22569 10625 22603 10659
rect 23489 10625 23523 10659
rect 25973 10625 26007 10659
rect 29285 10625 29319 10659
rect 30849 10625 30883 10659
rect 9597 10557 9631 10591
rect 11713 10557 11747 10591
rect 11989 10557 12023 10591
rect 13461 10557 13495 10591
rect 14013 10557 14047 10591
rect 18429 10557 18463 10591
rect 20177 10557 20211 10591
rect 24777 10557 24811 10591
rect 25789 10557 25823 10591
rect 10425 10489 10459 10523
rect 17233 10489 17267 10523
rect 6653 10421 6687 10455
rect 15761 10421 15795 10455
rect 23029 10421 23063 10455
rect 26157 10421 26191 10455
rect 30941 10421 30975 10455
rect 3433 10217 3467 10251
rect 16589 10217 16623 10251
rect 22477 10217 22511 10251
rect 25329 10217 25363 10251
rect 13645 10149 13679 10183
rect 20085 10149 20119 10183
rect 1685 10081 1719 10115
rect 3985 10081 4019 10115
rect 6837 10081 6871 10115
rect 7113 10081 7147 10115
rect 14657 10081 14691 10115
rect 15577 10081 15611 10115
rect 17325 10081 17359 10115
rect 18705 10081 18739 10115
rect 19534 10081 19568 10115
rect 23213 10081 23247 10115
rect 37749 10081 37783 10115
rect 6009 10013 6043 10047
rect 11897 10013 11931 10047
rect 16129 10013 16163 10047
rect 16313 10013 16347 10047
rect 18429 10013 18463 10047
rect 24777 10013 24811 10047
rect 25237 10013 25271 10047
rect 26065 10013 26099 10047
rect 37473 10013 37507 10047
rect 1961 9945 1995 9979
rect 4261 9945 4295 9979
rect 9137 9945 9171 9979
rect 12173 9945 12207 9979
rect 14749 9945 14783 9979
rect 17417 9945 17451 9979
rect 17969 9945 18003 9979
rect 19625 9945 19659 9979
rect 21189 9945 21223 9979
rect 21281 9945 21315 9979
rect 21833 9945 21867 9979
rect 22385 9945 22419 9979
rect 23305 9945 23339 9979
rect 23857 9945 23891 9979
rect 8585 9877 8619 9911
rect 10425 9877 10459 9911
rect 24593 9877 24627 9911
rect 25881 9877 25915 9911
rect 14381 9605 14415 9639
rect 17049 9605 17083 9639
rect 17601 9605 17635 9639
rect 18613 9605 18647 9639
rect 21465 9605 21499 9639
rect 22753 9605 22787 9639
rect 6745 9537 6779 9571
rect 9965 9537 9999 9571
rect 10701 9537 10735 9571
rect 15853 9537 15887 9571
rect 19625 9537 19659 9571
rect 22017 9537 22051 9571
rect 22661 9537 22695 9571
rect 23305 9537 23339 9571
rect 24501 9537 24535 9571
rect 25789 9537 25823 9571
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 6009 9469 6043 9503
rect 7481 9469 7515 9503
rect 7757 9469 7791 9503
rect 9505 9469 9539 9503
rect 11897 9469 11931 9503
rect 12173 9469 12207 9503
rect 13921 9469 13955 9503
rect 15117 9469 15151 9503
rect 16129 9469 16163 9503
rect 16957 9469 16991 9503
rect 18521 9469 18555 9503
rect 18797 9469 18831 9503
rect 19901 9469 19935 9503
rect 20821 9469 20855 9503
rect 21005 9469 21039 9503
rect 23397 9469 23431 9503
rect 24685 9469 24719 9503
rect 6561 9401 6595 9435
rect 25605 9401 25639 9435
rect 3341 9333 3375 9367
rect 22109 9333 22143 9367
rect 24869 9333 24903 9367
rect 2605 9129 2639 9163
rect 5641 9129 5675 9163
rect 9413 9129 9447 9163
rect 12357 9129 12391 9163
rect 20729 9129 20763 9163
rect 23857 9129 23891 9163
rect 24593 9129 24627 9163
rect 29837 9129 29871 9163
rect 3341 9061 3375 9095
rect 7941 9061 7975 9095
rect 4721 8993 4755 9027
rect 6469 8993 6503 9027
rect 10609 8993 10643 9027
rect 10885 8993 10919 9027
rect 14289 8993 14323 9027
rect 16037 8993 16071 9027
rect 17049 8993 17083 9027
rect 19533 9005 19567 9039
rect 19993 8993 20027 9027
rect 22569 8993 22603 9027
rect 1593 8925 1627 8959
rect 2789 8925 2823 8959
rect 3249 8925 3283 8959
rect 5549 8925 5583 8959
rect 6193 8925 6227 8959
rect 9321 8925 9355 8959
rect 10149 8925 10183 8959
rect 13277 8925 13311 8959
rect 16865 8925 16899 8959
rect 18705 8925 18739 8959
rect 20637 8925 20671 8959
rect 22477 8925 22511 8959
rect 23121 8925 23155 8959
rect 23765 8925 23799 8959
rect 24777 8925 24811 8959
rect 25237 8925 25271 8959
rect 29745 8925 29779 8959
rect 3985 8857 4019 8891
rect 13553 8857 13587 8891
rect 14565 8857 14599 8891
rect 18061 8857 18095 8891
rect 18153 8857 18187 8891
rect 19625 8857 19659 8891
rect 21373 8857 21407 8891
rect 21465 8857 21499 8891
rect 22017 8857 22051 8891
rect 1777 8789 1811 8823
rect 9965 8789 9999 8823
rect 17509 8789 17543 8823
rect 23213 8789 23247 8823
rect 25329 8789 25363 8823
rect 1777 8585 1811 8619
rect 5273 8585 5307 8619
rect 16221 8585 16255 8619
rect 17509 8585 17543 8619
rect 25145 8585 25179 8619
rect 38117 8585 38151 8619
rect 2697 8517 2731 8551
rect 6653 8517 6687 8551
rect 10149 8517 10183 8551
rect 14657 8517 14691 8551
rect 14749 8517 14783 8551
rect 18153 8517 18187 8551
rect 20085 8517 20119 8551
rect 21373 8517 21407 8551
rect 1961 8449 1995 8483
rect 5181 8449 5215 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 10057 8449 10091 8483
rect 10701 8449 10735 8483
rect 10977 8449 11011 8483
rect 11989 8449 12023 8483
rect 16129 8449 16163 8483
rect 16865 8449 16899 8483
rect 20637 8449 20671 8483
rect 21189 8449 21223 8483
rect 22017 8449 22051 8483
rect 24133 8449 24167 8483
rect 25053 8449 25087 8483
rect 25697 8449 25731 8483
rect 32965 8449 32999 8483
rect 38301 8449 38335 8483
rect 2421 8381 2455 8415
rect 4169 8381 4203 8415
rect 5917 8381 5951 8415
rect 7481 8381 7515 8415
rect 7757 8381 7791 8415
rect 9505 8381 9539 8415
rect 12265 8381 12299 8415
rect 14013 8381 14047 8415
rect 15669 8381 15703 8415
rect 17049 8381 17083 8415
rect 18061 8381 18095 8415
rect 18613 8381 18647 8415
rect 19993 8381 20027 8415
rect 23029 8381 23063 8415
rect 23213 8381 23247 8415
rect 24225 8381 24259 8415
rect 22109 8313 22143 8347
rect 23673 8313 23707 8347
rect 25789 8313 25823 8347
rect 33057 8313 33091 8347
rect 2973 8041 3007 8075
rect 23397 8041 23431 8075
rect 31401 8041 31435 8075
rect 7665 7973 7699 8007
rect 10885 7973 10919 8007
rect 16037 7973 16071 8007
rect 19717 7973 19751 8007
rect 24685 7973 24719 8007
rect 38117 7973 38151 8007
rect 1869 7905 1903 7939
rect 5089 7905 5123 7939
rect 9137 7905 9171 7939
rect 11621 7905 11655 7939
rect 13369 7905 13403 7939
rect 15209 7905 15243 7939
rect 16681 7905 16715 7939
rect 17601 7905 17635 7939
rect 20361 7905 20395 7939
rect 20821 7905 20855 7939
rect 21557 7905 21591 7939
rect 1593 7837 1627 7871
rect 2881 7837 2915 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 4721 7837 4755 7871
rect 5917 7837 5951 7871
rect 8401 7837 8435 7871
rect 11345 7837 11379 7871
rect 15853 7837 15887 7871
rect 18153 7837 18187 7871
rect 18429 7837 18463 7871
rect 22661 7837 22695 7871
rect 23305 7837 23339 7871
rect 24593 7837 24627 7871
rect 31309 7837 31343 7871
rect 35725 7837 35759 7871
rect 38301 7837 38335 7871
rect 6193 7769 6227 7803
rect 9413 7769 9447 7803
rect 14749 7769 14783 7803
rect 14841 7769 14875 7803
rect 16773 7769 16807 7803
rect 19533 7769 19567 7803
rect 20453 7769 20487 7803
rect 21649 7769 21683 7803
rect 22201 7769 22235 7803
rect 4077 7701 4111 7735
rect 5641 7701 5675 7735
rect 8493 7701 8527 7735
rect 35541 7701 35575 7735
rect 5273 7497 5307 7531
rect 22753 7497 22787 7531
rect 23397 7497 23431 7531
rect 25237 7497 25271 7531
rect 2513 7429 2547 7463
rect 7297 7429 7331 7463
rect 8585 7429 8619 7463
rect 14473 7429 14507 7463
rect 15301 7429 15335 7463
rect 17417 7429 17451 7463
rect 19441 7429 19475 7463
rect 20637 7429 20671 7463
rect 20729 7429 20763 7463
rect 22109 7429 22143 7463
rect 1777 7361 1811 7395
rect 2237 7361 2271 7395
rect 4537 7361 4571 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 6561 7361 6595 7395
rect 8309 7361 8343 7395
rect 10609 7361 10643 7395
rect 10701 7361 10735 7395
rect 14197 7361 14231 7395
rect 22017 7361 22051 7395
rect 22661 7361 22695 7395
rect 23305 7361 23339 7395
rect 24409 7361 24443 7395
rect 25421 7361 25455 7395
rect 3985 7293 4019 7327
rect 5917 7293 5951 7327
rect 11897 7293 11931 7327
rect 12173 7293 12207 7327
rect 15209 7293 15243 7327
rect 17325 7293 17359 7327
rect 17785 7293 17819 7327
rect 19349 7293 19383 7327
rect 20913 7293 20947 7327
rect 23949 7293 23983 7327
rect 24869 7293 24903 7327
rect 4629 7225 4663 7259
rect 15761 7225 15795 7259
rect 19901 7225 19935 7259
rect 1593 7157 1627 7191
rect 10057 7157 10091 7191
rect 13645 7157 13679 7191
rect 24501 7157 24535 7191
rect 1856 6953 1890 6987
rect 6174 6953 6208 6987
rect 7665 6953 7699 6987
rect 8493 6885 8527 6919
rect 3341 6817 3375 6851
rect 13553 6817 13587 6851
rect 14381 6817 14415 6851
rect 15025 6817 15059 6851
rect 15669 6817 15703 6851
rect 16681 6817 16715 6851
rect 17325 6817 17359 6851
rect 19533 6817 19567 6851
rect 21373 6817 21407 6851
rect 22385 6817 22419 6851
rect 23397 6817 23431 6851
rect 1593 6749 1627 6783
rect 4261 6749 4295 6783
rect 5917 6749 5951 6783
rect 8393 6751 8427 6785
rect 9413 6749 9447 6783
rect 10057 6749 10091 6783
rect 12357 6749 12391 6783
rect 13277 6749 13311 6783
rect 14289 6749 14323 6783
rect 20177 6749 20211 6783
rect 21189 6749 21223 6783
rect 22293 6749 22327 6783
rect 23581 6749 23615 6783
rect 24593 6749 24627 6783
rect 4997 6681 5031 6715
rect 10333 6681 10367 6715
rect 12633 6681 12667 6715
rect 15117 6681 15151 6715
rect 16773 6681 16807 6715
rect 18153 6681 18187 6715
rect 18245 6681 18279 6715
rect 18797 6681 18831 6715
rect 19625 6681 19659 6715
rect 9505 6613 9539 6647
rect 11805 6613 11839 6647
rect 21833 6613 21867 6647
rect 24041 6613 24075 6647
rect 24685 6613 24719 6647
rect 21005 6409 21039 6443
rect 22753 6409 22787 6443
rect 27169 6409 27203 6443
rect 32413 6409 32447 6443
rect 38117 6409 38151 6443
rect 7205 6341 7239 6375
rect 9413 6341 9447 6375
rect 14197 6341 14231 6375
rect 15117 6341 15151 6375
rect 15761 6341 15795 6375
rect 17693 6341 17727 6375
rect 18797 6341 18831 6375
rect 19901 6341 19935 6375
rect 23397 6341 23431 6375
rect 24685 6341 24719 6375
rect 1961 6273 1995 6307
rect 2973 6273 3007 6307
rect 3065 6273 3099 6307
rect 3801 6273 3835 6307
rect 4261 6273 4295 6307
rect 6929 6273 6963 6307
rect 9137 6273 9171 6307
rect 16313 6273 16347 6307
rect 16865 6273 16899 6307
rect 18245 6273 18279 6307
rect 18705 6273 18739 6307
rect 20453 6273 20487 6307
rect 20913 6273 20947 6307
rect 22017 6273 22051 6307
rect 22109 6273 22143 6307
rect 22661 6273 22695 6307
rect 23305 6273 23339 6307
rect 23949 6273 23983 6307
rect 24593 6273 24627 6307
rect 25329 6273 25363 6307
rect 26157 6273 26191 6307
rect 27353 6273 27387 6307
rect 32321 6273 32355 6307
rect 38301 6273 38335 6307
rect 4537 6205 4571 6239
rect 10885 6205 10919 6239
rect 11713 6205 11747 6239
rect 11989 6205 12023 6239
rect 14105 6205 14139 6239
rect 15669 6205 15703 6239
rect 16957 6205 16991 6239
rect 17601 6205 17635 6239
rect 19809 6205 19843 6239
rect 3617 6137 3651 6171
rect 24041 6137 24075 6171
rect 1777 6069 1811 6103
rect 6009 6069 6043 6103
rect 8677 6069 8711 6103
rect 13461 6069 13495 6103
rect 25421 6069 25455 6103
rect 25973 6069 26007 6103
rect 5917 5865 5951 5899
rect 8585 5865 8619 5899
rect 23857 5865 23891 5899
rect 24869 5865 24903 5899
rect 26433 5865 26467 5899
rect 10609 5797 10643 5831
rect 13001 5797 13035 5831
rect 19809 5797 19843 5831
rect 21925 5797 21959 5831
rect 23213 5797 23247 5831
rect 24501 5797 24535 5831
rect 1685 5729 1719 5763
rect 4169 5729 4203 5763
rect 7113 5729 7147 5763
rect 9873 5729 9907 5763
rect 11253 5729 11287 5763
rect 11529 5729 11563 5763
rect 14289 5729 14323 5763
rect 18245 5729 18279 5763
rect 20637 5729 20671 5763
rect 21281 5729 21315 5763
rect 6837 5661 6871 5695
rect 10517 5661 10551 5695
rect 13553 5661 13587 5695
rect 16681 5661 16715 5695
rect 19441 5661 19475 5695
rect 19625 5661 19659 5695
rect 20545 5661 20579 5695
rect 21189 5661 21223 5695
rect 21833 5661 21867 5695
rect 22477 5661 22511 5695
rect 23121 5661 23155 5695
rect 23765 5661 23799 5695
rect 24409 5661 24443 5695
rect 25421 5661 25455 5695
rect 26617 5661 26651 5695
rect 1961 5593 1995 5627
rect 4445 5593 4479 5627
rect 9137 5593 9171 5627
rect 14565 5593 14599 5627
rect 17417 5593 17451 5627
rect 17509 5593 17543 5627
rect 3433 5525 3467 5559
rect 13645 5525 13679 5559
rect 16037 5525 16071 5559
rect 16681 5525 16715 5559
rect 22569 5525 22603 5559
rect 25237 5525 25271 5559
rect 24685 5321 24719 5355
rect 4537 5253 4571 5287
rect 13921 5253 13955 5287
rect 14657 5253 14691 5287
rect 15761 5253 15795 5287
rect 17325 5253 17359 5287
rect 18521 5253 18555 5287
rect 19073 5253 19107 5287
rect 19809 5253 19843 5287
rect 4261 5185 4295 5219
rect 6561 5185 6595 5219
rect 7205 5185 7239 5219
rect 16313 5185 16347 5219
rect 21089 5175 21123 5209
rect 22661 5185 22695 5219
rect 23305 5185 23339 5219
rect 23949 5185 23983 5219
rect 24593 5185 24627 5219
rect 25421 5185 25455 5219
rect 38025 5185 38059 5219
rect 2053 5117 2087 5151
rect 2329 5117 2363 5151
rect 3801 5117 3835 5151
rect 7481 5117 7515 5151
rect 9413 5117 9447 5151
rect 9689 5117 9723 5151
rect 11713 5117 11747 5151
rect 11989 5117 12023 5151
rect 15669 5117 15703 5151
rect 17233 5117 17267 5151
rect 18429 5117 18463 5151
rect 19717 5117 19751 5151
rect 20361 5117 20395 5151
rect 22017 5117 22051 5151
rect 22753 5117 22787 5151
rect 6009 5049 6043 5083
rect 11161 5049 11195 5083
rect 17785 5049 17819 5083
rect 23397 5049 23431 5083
rect 6653 4981 6687 5015
rect 8953 4981 8987 5015
rect 13461 4981 13495 5015
rect 21189 4981 21223 5015
rect 24041 4981 24075 5015
rect 25237 4981 25271 5015
rect 38209 4981 38243 5015
rect 1856 4777 1890 4811
rect 7849 4777 7883 4811
rect 11332 4777 11366 4811
rect 12817 4777 12851 4811
rect 13645 4777 13679 4811
rect 18521 4777 18555 4811
rect 19809 4777 19843 4811
rect 20545 4777 20579 4811
rect 21281 4777 21315 4811
rect 23213 4777 23247 4811
rect 28181 4777 28215 4811
rect 38117 4777 38151 4811
rect 3341 4709 3375 4743
rect 6653 4709 6687 4743
rect 25881 4709 25915 4743
rect 1593 4641 1627 4675
rect 4905 4641 4939 4675
rect 8493 4641 8527 4675
rect 14289 4641 14323 4675
rect 16957 4641 16991 4675
rect 17969 4641 18003 4675
rect 19441 4641 19475 4675
rect 19625 4641 19659 4675
rect 31493 4641 31527 4675
rect 4445 4573 4479 4607
rect 7757 4573 7791 4607
rect 8401 4573 8435 4607
rect 9689 4573 9723 4607
rect 10517 4573 10551 4607
rect 11069 4573 11103 4607
rect 13553 4573 13587 4607
rect 18429 4573 18463 4607
rect 20729 4573 20763 4607
rect 21189 4573 21223 4607
rect 21833 4573 21867 4607
rect 22477 4573 22511 4607
rect 23121 4573 23155 4607
rect 23765 4573 23799 4607
rect 23857 4573 23891 4607
rect 24685 4573 24719 4607
rect 25237 4573 25271 4607
rect 25329 4573 25363 4607
rect 26065 4573 26099 4607
rect 26341 4573 26375 4607
rect 28089 4573 28123 4607
rect 30941 4573 30975 4607
rect 31401 4573 31435 4607
rect 38301 4573 38335 4607
rect 5181 4505 5215 4539
rect 14565 4505 14599 4539
rect 17042 4505 17076 4539
rect 22569 4505 22603 4539
rect 25421 4505 25455 4539
rect 4261 4437 4295 4471
rect 16037 4437 16071 4471
rect 21925 4437 21959 4471
rect 25053 4437 25087 4471
rect 30757 4437 30791 4471
rect 19901 4233 19935 4267
rect 20361 4233 20395 4267
rect 21097 4233 21131 4267
rect 22753 4233 22787 4267
rect 25329 4233 25363 4267
rect 3433 4165 3467 4199
rect 14473 4165 14507 4199
rect 17325 4165 17359 4199
rect 38117 4165 38151 4199
rect 1593 4097 1627 4131
rect 2513 4097 2547 4131
rect 3157 4097 3191 4131
rect 5825 4097 5859 4131
rect 5917 4097 5951 4131
rect 6653 4097 6687 4131
rect 14197 4097 14231 4131
rect 20545 4097 20579 4131
rect 21005 4097 21039 4131
rect 22017 4097 22051 4131
rect 22661 4097 22695 4131
rect 23305 4097 23339 4131
rect 23949 4097 23983 4131
rect 24593 4097 24627 4131
rect 25237 4097 25271 4131
rect 27353 4097 27387 4131
rect 4905 4029 4939 4063
rect 6929 4029 6963 4063
rect 9321 4029 9355 4063
rect 11713 4029 11747 4063
rect 11989 4029 12023 4063
rect 13737 4029 13771 4063
rect 17233 4029 17267 4063
rect 18245 4029 18279 4063
rect 19257 4029 19291 4063
rect 19441 4029 19475 4063
rect 1777 3961 1811 3995
rect 11069 3961 11103 3995
rect 22109 3961 22143 3995
rect 26065 3961 26099 3995
rect 2605 3893 2639 3927
rect 8401 3893 8435 3927
rect 9584 3893 9618 3927
rect 15945 3893 15979 3927
rect 23397 3893 23431 3927
rect 24041 3893 24075 3927
rect 24685 3893 24719 3927
rect 27169 3893 27203 3927
rect 38209 3893 38243 3927
rect 2237 3689 2271 3723
rect 8493 3689 8527 3723
rect 9781 3689 9815 3723
rect 10596 3689 10630 3723
rect 13001 3689 13035 3723
rect 13645 3689 13679 3723
rect 20177 3689 20211 3723
rect 25973 3689 26007 3723
rect 3341 3621 3375 3655
rect 7205 3621 7239 3655
rect 21465 3621 21499 3655
rect 22109 3621 22143 3655
rect 37565 3621 37599 3655
rect 10333 3553 10367 3587
rect 12357 3553 12391 3587
rect 15669 3553 15703 3587
rect 19533 3553 19567 3587
rect 20821 3553 20855 3587
rect 1593 3485 1627 3519
rect 2605 3485 2639 3519
rect 3249 3485 3283 3519
rect 4537 3485 4571 3519
rect 6561 3485 6595 3519
rect 7113 3485 7147 3519
rect 7757 3485 7791 3519
rect 8401 3485 8435 3519
rect 9689 3485 9723 3519
rect 12909 3485 12943 3519
rect 13553 3485 13587 3519
rect 16773 3485 16807 3519
rect 16865 3485 16899 3519
rect 18429 3485 18463 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 20729 3485 20763 3519
rect 21373 3485 21407 3519
rect 22017 3485 22051 3519
rect 22661 3485 22695 3519
rect 22753 3485 22787 3519
rect 23489 3485 23523 3519
rect 24593 3485 24627 3519
rect 25237 3485 25271 3519
rect 25881 3485 25915 3519
rect 26525 3485 26559 3519
rect 27353 3485 27387 3519
rect 27997 3485 28031 3519
rect 38025 3485 38059 3519
rect 4813 3417 4847 3451
rect 14473 3417 14507 3451
rect 14565 3417 14599 3451
rect 15117 3417 15151 3451
rect 15761 3417 15795 3451
rect 16313 3417 16347 3451
rect 17785 3417 17819 3451
rect 17877 3417 17911 3451
rect 37381 3417 37415 3451
rect 1777 3349 1811 3383
rect 2697 3349 2731 3383
rect 7849 3349 7883 3383
rect 23305 3349 23339 3383
rect 24685 3349 24719 3383
rect 25329 3349 25363 3383
rect 26617 3349 26651 3383
rect 27169 3349 27203 3383
rect 27813 3349 27847 3383
rect 38209 3349 38243 3383
rect 3341 3145 3375 3179
rect 5273 3145 5307 3179
rect 6837 3145 6871 3179
rect 8769 3145 8803 3179
rect 10425 3145 10459 3179
rect 11069 3145 11103 3179
rect 14749 3145 14783 3179
rect 15393 3145 15427 3179
rect 16037 3145 16071 3179
rect 18429 3145 18463 3179
rect 19073 3145 19107 3179
rect 19717 3145 19751 3179
rect 27813 3145 27847 3179
rect 36737 3145 36771 3179
rect 4629 3077 4663 3111
rect 5917 3077 5951 3111
rect 17233 3077 17267 3111
rect 17325 3077 17359 3111
rect 24869 3077 24903 3111
rect 25513 3077 25547 3111
rect 1593 3009 1627 3043
rect 2329 3009 2363 3043
rect 3249 3009 3283 3043
rect 3893 3009 3927 3043
rect 4537 3009 4571 3043
rect 5181 3009 5215 3043
rect 5825 3009 5859 3043
rect 6753 3015 6787 3049
rect 7389 3009 7423 3043
rect 8033 3009 8067 3043
rect 8677 3009 8711 3043
rect 9321 3009 9355 3043
rect 10333 3009 10367 3043
rect 10977 3009 11011 3043
rect 11805 3009 11839 3043
rect 14013 3009 14047 3043
rect 14657 3009 14691 3043
rect 15309 3009 15343 3043
rect 15945 3009 15979 3043
rect 18337 3009 18371 3043
rect 18981 3009 19015 3043
rect 19633 3007 19667 3041
rect 20269 3009 20303 3043
rect 20361 3009 20395 3043
rect 21097 3009 21131 3043
rect 22201 3009 22235 3043
rect 22661 3009 22695 3043
rect 23489 3009 23523 3043
rect 23949 3009 23983 3043
rect 24777 3009 24811 3043
rect 25421 3009 25455 3043
rect 26249 3009 26283 3043
rect 27169 3009 27203 3043
rect 27997 3009 28031 3043
rect 36921 3009 36955 3043
rect 37749 3009 37783 3043
rect 3985 2941 4019 2975
rect 7481 2941 7515 2975
rect 9413 2941 9447 2975
rect 12081 2941 12115 2975
rect 13553 2941 13587 2975
rect 17877 2941 17911 2975
rect 24041 2941 24075 2975
rect 37473 2941 37507 2975
rect 2513 2873 2547 2907
rect 22017 2873 22051 2907
rect 1777 2805 1811 2839
rect 8125 2805 8159 2839
rect 14105 2805 14139 2839
rect 20913 2805 20947 2839
rect 22753 2805 22787 2839
rect 23305 2805 23339 2839
rect 26065 2805 26099 2839
rect 27261 2805 27295 2839
rect 7849 2601 7883 2635
rect 10517 2601 10551 2635
rect 13737 2601 13771 2635
rect 14841 2601 14875 2635
rect 16129 2601 16163 2635
rect 16957 2601 16991 2635
rect 17601 2601 17635 2635
rect 20177 2601 20211 2635
rect 22017 2601 22051 2635
rect 24593 2601 24627 2635
rect 27169 2601 27203 2635
rect 28457 2601 28491 2635
rect 30481 2601 30515 2635
rect 32321 2601 32355 2635
rect 33149 2601 33183 2635
rect 20729 2533 20763 2567
rect 4261 2465 4295 2499
rect 9413 2465 9447 2499
rect 11989 2465 12023 2499
rect 12265 2465 12299 2499
rect 2053 2397 2087 2431
rect 3157 2397 3191 2431
rect 3985 2397 4019 2431
rect 5273 2397 5307 2431
rect 6561 2397 6595 2431
rect 7757 2397 7791 2431
rect 8401 2397 8435 2431
rect 9137 2397 9171 2431
rect 10425 2397 10459 2431
rect 14749 2397 14783 2431
rect 15393 2397 15427 2431
rect 16037 2397 16071 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 18153 2397 18187 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 20913 2397 20947 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 25973 2397 26007 2431
rect 27353 2397 27387 2431
rect 28641 2397 28675 2431
rect 29745 2397 29779 2431
rect 30665 2397 30699 2431
rect 32505 2397 32539 2431
rect 33701 2397 33735 2431
rect 34897 2397 34931 2431
rect 36185 2397 36219 2431
rect 37473 2397 37507 2431
rect 37749 2397 37783 2431
rect 33057 2329 33091 2363
rect 2237 2261 2271 2295
rect 3341 2261 3375 2295
rect 5457 2261 5491 2295
rect 6745 2261 6779 2295
rect 8493 2261 8527 2295
rect 15485 2261 15519 2295
rect 18337 2261 18371 2295
rect 19533 2261 19567 2295
rect 22845 2261 22879 2295
rect 23397 2261 23431 2295
rect 25421 2261 25455 2295
rect 26157 2261 26191 2295
rect 29929 2261 29963 2295
rect 33885 2261 33919 2295
rect 35081 2261 35115 2295
rect 36369 2261 36403 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1578 37312 1584 37324
rect 1539 37284 1584 37312
rect 1578 37272 1584 37284
rect 1636 37272 1642 37324
rect 9493 37315 9551 37321
rect 4540 37284 4936 37312
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37213 1915 37247
rect 2866 37244 2872 37256
rect 2827 37216 2872 37244
rect 1857 37207 1915 37213
rect 1872 37176 1900 37207
rect 2866 37204 2872 37216
rect 2924 37204 2930 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 4157 37247 4215 37253
rect 4157 37244 4169 37247
rect 3292 37216 4169 37244
rect 3292 37204 3298 37216
rect 4157 37213 4169 37216
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4540 37176 4568 37284
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4801 37247 4859 37253
rect 4801 37244 4813 37247
rect 4672 37216 4813 37244
rect 4672 37204 4678 37216
rect 4801 37213 4813 37216
rect 4847 37213 4859 37247
rect 4908 37244 4936 37284
rect 9493 37281 9505 37315
rect 9539 37312 9551 37315
rect 9539 37284 9812 37312
rect 9539 37281 9551 37284
rect 9493 37275 9551 37281
rect 9784 37256 9812 37284
rect 10962 37272 10968 37324
rect 11020 37312 11026 37324
rect 11701 37315 11759 37321
rect 11701 37312 11713 37315
rect 11020 37284 11713 37312
rect 11020 37272 11026 37284
rect 11701 37281 11713 37284
rect 11747 37281 11759 37315
rect 11701 37275 11759 37281
rect 21266 37272 21272 37324
rect 21324 37312 21330 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 21324 37284 22017 37312
rect 21324 37272 21330 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 30926 37312 30932 37324
rect 30887 37284 30932 37312
rect 22005 37275 22063 37281
rect 30926 37272 30932 37284
rect 30984 37272 30990 37324
rect 34146 37272 34152 37324
rect 34204 37312 34210 37324
rect 34885 37315 34943 37321
rect 34885 37312 34897 37315
rect 34204 37284 34897 37312
rect 34204 37272 34210 37284
rect 34885 37281 34897 37284
rect 34931 37281 34943 37315
rect 34885 37275 34943 37281
rect 37461 37315 37519 37321
rect 37461 37281 37473 37315
rect 37507 37312 37519 37315
rect 38654 37312 38660 37324
rect 37507 37284 38660 37312
rect 37507 37281 37519 37284
rect 37461 37275 37519 37281
rect 38654 37272 38660 37284
rect 38712 37272 38718 37324
rect 5534 37244 5540 37256
rect 4908 37216 5540 37244
rect 4801 37207 4859 37213
rect 5534 37204 5540 37216
rect 5592 37204 5598 37256
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 5997 37247 6055 37253
rect 5997 37244 6009 37247
rect 5868 37216 6009 37244
rect 5868 37204 5874 37216
rect 5997 37213 6009 37216
rect 6043 37213 6055 37247
rect 5997 37207 6055 37213
rect 6454 37204 6460 37256
rect 6512 37244 6518 37256
rect 6733 37247 6791 37253
rect 6733 37244 6745 37247
rect 6512 37216 6745 37244
rect 6512 37204 6518 37216
rect 6733 37213 6745 37216
rect 6779 37213 6791 37247
rect 7834 37244 7840 37256
rect 7795 37216 7840 37244
rect 6733 37207 6791 37213
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 9766 37244 9772 37256
rect 9727 37216 9772 37244
rect 9766 37204 9772 37216
rect 9824 37204 9830 37256
rect 11790 37204 11796 37256
rect 11848 37244 11854 37256
rect 11977 37247 12035 37253
rect 11977 37244 11989 37247
rect 11848 37216 11989 37244
rect 11848 37204 11854 37216
rect 11977 37213 11989 37216
rect 12023 37213 12035 37247
rect 11977 37207 12035 37213
rect 12434 37204 12440 37256
rect 12492 37244 12498 37256
rect 13173 37247 13231 37253
rect 13173 37244 13185 37247
rect 12492 37216 13185 37244
rect 12492 37204 12498 37216
rect 13173 37213 13185 37216
rect 13219 37213 13231 37247
rect 14274 37244 14280 37256
rect 14235 37216 14280 37244
rect 13173 37207 13231 37213
rect 14274 37204 14280 37216
rect 14332 37204 14338 37256
rect 15470 37204 15476 37256
rect 15528 37244 15534 37256
rect 15749 37247 15807 37253
rect 15749 37244 15761 37247
rect 15528 37216 15761 37244
rect 15528 37204 15534 37216
rect 15749 37213 15761 37216
rect 15795 37213 15807 37247
rect 17494 37244 17500 37256
rect 17455 37216 17500 37244
rect 15749 37207 15807 37213
rect 17494 37204 17500 37216
rect 17552 37204 17558 37256
rect 19426 37204 19432 37256
rect 19484 37244 19490 37256
rect 19613 37247 19671 37253
rect 19613 37244 19625 37247
rect 19484 37216 19625 37244
rect 19484 37204 19490 37216
rect 19613 37213 19625 37216
rect 19659 37213 19671 37247
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 19613 37207 19671 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 22281 37247 22339 37253
rect 22281 37213 22293 37247
rect 22327 37213 22339 37247
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 22281 37207 22339 37213
rect 9398 37176 9404 37188
rect 1872 37148 4568 37176
rect 4632 37148 9404 37176
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 3053 37111 3111 37117
rect 3053 37108 3065 37111
rect 2832 37080 3065 37108
rect 2832 37068 2838 37080
rect 3053 37077 3065 37080
rect 3099 37077 3111 37111
rect 3970 37108 3976 37120
rect 3931 37080 3976 37108
rect 3053 37071 3111 37077
rect 3970 37068 3976 37080
rect 4028 37068 4034 37120
rect 4632 37117 4660 37148
rect 9398 37136 9404 37148
rect 9456 37136 9462 37188
rect 18782 37136 18788 37188
rect 18840 37176 18846 37188
rect 22296 37176 22324 37207
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 25130 37204 25136 37256
rect 25188 37244 25194 37256
rect 25501 37247 25559 37253
rect 25501 37244 25513 37247
rect 25188 37216 25513 37244
rect 25188 37204 25194 37216
rect 25501 37213 25513 37216
rect 25547 37213 25559 37247
rect 25501 37207 25559 37213
rect 26418 37204 26424 37256
rect 26476 37244 26482 37256
rect 27341 37247 27399 37253
rect 27341 37244 27353 37247
rect 26476 37216 27353 37244
rect 26476 37204 26482 37216
rect 27341 37213 27353 37216
rect 27387 37213 27399 37247
rect 27798 37244 27804 37256
rect 27759 37216 27804 37244
rect 27341 37207 27399 37213
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 28350 37204 28356 37256
rect 28408 37244 28414 37256
rect 28721 37247 28779 37253
rect 28721 37244 28733 37247
rect 28408 37216 28733 37244
rect 28408 37204 28414 37216
rect 28721 37213 28733 37216
rect 28767 37213 28779 37247
rect 28721 37207 28779 37213
rect 29638 37204 29644 37256
rect 29696 37244 29702 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29696 37216 29929 37244
rect 29696 37204 29702 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 31205 37247 31263 37253
rect 31205 37213 31217 37247
rect 31251 37213 31263 37247
rect 32306 37244 32312 37256
rect 32267 37216 32312 37244
rect 31205 37207 31263 37213
rect 18840 37148 22324 37176
rect 18840 37136 18846 37148
rect 22370 37136 22376 37188
rect 22428 37176 22434 37188
rect 31220 37176 31248 37207
rect 32306 37204 32312 37216
rect 32364 37204 32370 37256
rect 32858 37204 32864 37256
rect 32916 37244 32922 37256
rect 33229 37247 33287 37253
rect 33229 37244 33241 37247
rect 32916 37216 33241 37244
rect 32916 37204 32922 37216
rect 33229 37213 33241 37216
rect 33275 37213 33287 37247
rect 33229 37207 33287 37213
rect 35161 37247 35219 37253
rect 35161 37213 35173 37247
rect 35207 37244 35219 37247
rect 35434 37244 35440 37256
rect 35207 37216 35440 37244
rect 35207 37213 35219 37216
rect 35161 37207 35219 37213
rect 35434 37204 35440 37216
rect 35492 37204 35498 37256
rect 35986 37204 35992 37256
rect 36044 37244 36050 37256
rect 36173 37247 36231 37253
rect 36173 37244 36185 37247
rect 36044 37216 36185 37244
rect 36044 37204 36050 37216
rect 36173 37213 36185 37216
rect 36219 37213 36231 37247
rect 36173 37207 36231 37213
rect 37737 37247 37795 37253
rect 37737 37213 37749 37247
rect 37783 37213 37795 37247
rect 37737 37207 37795 37213
rect 22428 37148 31248 37176
rect 22428 37136 22434 37148
rect 31294 37136 31300 37188
rect 31352 37176 31358 37188
rect 37752 37176 37780 37207
rect 31352 37148 37780 37176
rect 31352 37136 31358 37148
rect 4617 37111 4675 37117
rect 4617 37077 4629 37111
rect 4663 37077 4675 37111
rect 5810 37108 5816 37120
rect 5771 37080 5816 37108
rect 4617 37071 4675 37077
rect 5810 37068 5816 37080
rect 5868 37068 5874 37120
rect 6546 37108 6552 37120
rect 6507 37080 6552 37108
rect 6546 37068 6552 37080
rect 6604 37068 6610 37120
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7800 37080 8033 37108
rect 7800 37068 7806 37080
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 8021 37071 8079 37077
rect 9674 37068 9680 37120
rect 9732 37108 9738 37120
rect 9953 37111 10011 37117
rect 9953 37108 9965 37111
rect 9732 37080 9965 37108
rect 9732 37068 9738 37080
rect 9953 37077 9965 37080
rect 9999 37077 10011 37111
rect 9953 37071 10011 37077
rect 12342 37068 12348 37120
rect 12400 37108 12406 37120
rect 12989 37111 13047 37117
rect 12989 37108 13001 37111
rect 12400 37080 13001 37108
rect 12400 37068 12406 37080
rect 12989 37077 13001 37080
rect 13035 37077 13047 37111
rect 12989 37071 13047 37077
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 13596 37080 14473 37108
rect 13596 37068 13602 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 15562 37108 15568 37120
rect 15523 37080 15568 37108
rect 14461 37071 14519 37077
rect 15562 37068 15568 37080
rect 15620 37068 15626 37120
rect 17402 37068 17408 37120
rect 17460 37108 17466 37120
rect 17681 37111 17739 37117
rect 17681 37108 17693 37111
rect 17460 37080 17693 37108
rect 17460 37068 17466 37080
rect 17681 37077 17693 37080
rect 17727 37077 17739 37111
rect 17681 37071 17739 37077
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19429 37111 19487 37117
rect 19429 37108 19441 37111
rect 19392 37080 19441 37108
rect 19392 37068 19398 37080
rect 19429 37077 19441 37080
rect 19475 37077 19487 37111
rect 19429 37071 19487 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 25314 37108 25320 37120
rect 25275 37080 25320 37108
rect 24765 37071 24823 37077
rect 25314 37068 25320 37080
rect 25372 37068 25378 37120
rect 27154 37108 27160 37120
rect 27115 37080 27160 37108
rect 27154 37068 27160 37080
rect 27212 37068 27218 37120
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 27764 37080 27997 37108
rect 27764 37068 27770 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 28534 37108 28540 37120
rect 28495 37080 28540 37108
rect 27985 37071 28043 37077
rect 28534 37068 28540 37080
rect 28592 37068 28598 37120
rect 28626 37068 28632 37120
rect 28684 37108 28690 37120
rect 29733 37111 29791 37117
rect 29733 37108 29745 37111
rect 28684 37080 29745 37108
rect 28684 37068 28690 37080
rect 29733 37077 29745 37080
rect 29779 37077 29791 37111
rect 29733 37071 29791 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 33042 37108 33048 37120
rect 33003 37080 33048 37108
rect 32493 37071 32551 37077
rect 33042 37068 33048 37080
rect 33100 37068 33106 37120
rect 35526 37068 35532 37120
rect 35584 37108 35590 37120
rect 36357 37111 36415 37117
rect 36357 37108 36369 37111
rect 35584 37080 36369 37108
rect 35584 37068 35590 37080
rect 36357 37077 36369 37080
rect 36403 37077 36415 37111
rect 36357 37071 36415 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 9030 36864 9036 36916
rect 9088 36904 9094 36916
rect 9309 36907 9367 36913
rect 9309 36904 9321 36907
rect 9088 36876 9321 36904
rect 9088 36864 9094 36876
rect 9309 36873 9321 36876
rect 9355 36873 9367 36907
rect 9309 36867 9367 36873
rect 13173 36907 13231 36913
rect 13173 36873 13185 36907
rect 13219 36904 13231 36907
rect 14274 36904 14280 36916
rect 13219 36876 14280 36904
rect 13219 36873 13231 36876
rect 13173 36867 13231 36873
rect 14274 36864 14280 36876
rect 14332 36864 14338 36916
rect 16758 36864 16764 36916
rect 16816 36904 16822 36916
rect 17037 36907 17095 36913
rect 17037 36904 17049 36907
rect 16816 36876 17049 36904
rect 16816 36864 16822 36876
rect 17037 36873 17049 36876
rect 17083 36873 17095 36907
rect 17037 36867 17095 36873
rect 22094 36864 22100 36916
rect 22152 36904 22158 36916
rect 22189 36907 22247 36913
rect 22189 36904 22201 36907
rect 22152 36876 22201 36904
rect 22152 36864 22158 36876
rect 22189 36873 22201 36876
rect 22235 36873 22247 36907
rect 22189 36867 22247 36873
rect 26053 36907 26111 36913
rect 26053 36873 26065 36907
rect 26099 36904 26111 36907
rect 27798 36904 27804 36916
rect 26099 36876 27804 36904
rect 26099 36873 26111 36876
rect 26053 36867 26111 36873
rect 27798 36864 27804 36876
rect 27856 36864 27862 36916
rect 36817 36907 36875 36913
rect 36817 36873 36829 36907
rect 36863 36904 36875 36907
rect 39298 36904 39304 36916
rect 36863 36876 39304 36904
rect 36863 36873 36875 36876
rect 36817 36867 36875 36873
rect 39298 36864 39304 36876
rect 39356 36864 39362 36916
rect 1302 36796 1308 36848
rect 1360 36836 1366 36848
rect 1360 36808 3096 36836
rect 1360 36796 1366 36808
rect 14 36728 20 36780
rect 72 36768 78 36780
rect 3068 36777 3096 36808
rect 14182 36796 14188 36848
rect 14240 36836 14246 36848
rect 14240 36808 14504 36836
rect 14240 36796 14246 36808
rect 1581 36771 1639 36777
rect 1581 36768 1593 36771
rect 72 36740 1593 36768
rect 72 36728 78 36740
rect 1581 36737 1593 36740
rect 1627 36737 1639 36771
rect 1581 36731 1639 36737
rect 3053 36771 3111 36777
rect 3053 36737 3065 36771
rect 3099 36737 3111 36771
rect 3053 36731 3111 36737
rect 8849 36771 8907 36777
rect 8849 36737 8861 36771
rect 8895 36768 8907 36771
rect 9122 36768 9128 36780
rect 8895 36740 9128 36768
rect 8895 36737 8907 36740
rect 8849 36731 8907 36737
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 13357 36771 13415 36777
rect 13357 36737 13369 36771
rect 13403 36768 13415 36771
rect 13538 36768 13544 36780
rect 13403 36740 13544 36768
rect 13403 36737 13415 36740
rect 13357 36731 13415 36737
rect 13538 36728 13544 36740
rect 13596 36768 13602 36780
rect 14476 36777 14504 36808
rect 19150 36796 19156 36848
rect 19208 36836 19214 36848
rect 22370 36836 22376 36848
rect 19208 36808 22376 36836
rect 19208 36796 19214 36808
rect 22370 36796 22376 36808
rect 22428 36796 22434 36848
rect 36078 36836 36084 36848
rect 35866 36808 36084 36836
rect 14461 36771 14519 36777
rect 13596 36740 14320 36768
rect 13596 36728 13602 36740
rect 1854 36700 1860 36712
rect 1815 36672 1860 36700
rect 1854 36660 1860 36672
rect 1912 36660 1918 36712
rect 14292 36641 14320 36740
rect 14461 36737 14473 36771
rect 14507 36737 14519 36771
rect 14461 36731 14519 36737
rect 15378 36728 15384 36780
rect 15436 36768 15442 36780
rect 16853 36771 16911 36777
rect 16853 36768 16865 36771
rect 15436 36740 16865 36768
rect 15436 36728 15442 36740
rect 16853 36737 16865 36740
rect 16899 36737 16911 36771
rect 16853 36731 16911 36737
rect 18046 36728 18052 36780
rect 18104 36768 18110 36780
rect 22005 36771 22063 36777
rect 22005 36768 22017 36771
rect 18104 36740 22017 36768
rect 18104 36728 18110 36740
rect 22005 36737 22017 36740
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 23198 36728 23204 36780
rect 23256 36768 23262 36780
rect 23293 36771 23351 36777
rect 23293 36768 23305 36771
rect 23256 36740 23305 36768
rect 23256 36728 23262 36740
rect 23293 36737 23305 36740
rect 23339 36737 23351 36771
rect 23293 36731 23351 36737
rect 26234 36728 26240 36780
rect 26292 36768 26298 36780
rect 31294 36768 31300 36780
rect 26292 36740 31300 36768
rect 26292 36728 26298 36740
rect 31294 36728 31300 36740
rect 31352 36728 31358 36780
rect 35529 36771 35587 36777
rect 35529 36737 35541 36771
rect 35575 36768 35587 36771
rect 35866 36768 35894 36808
rect 36078 36796 36084 36808
rect 36136 36796 36142 36848
rect 38102 36836 38108 36848
rect 38063 36808 38108 36836
rect 38102 36796 38108 36808
rect 38160 36796 38166 36848
rect 36170 36768 36176 36780
rect 35575 36740 35894 36768
rect 36131 36740 36176 36768
rect 35575 36737 35587 36740
rect 35529 36731 35587 36737
rect 36170 36728 36176 36740
rect 36228 36728 36234 36780
rect 36633 36771 36691 36777
rect 36633 36737 36645 36771
rect 36679 36737 36691 36771
rect 36633 36731 36691 36737
rect 20622 36660 20628 36712
rect 20680 36700 20686 36712
rect 23569 36703 23627 36709
rect 23569 36700 23581 36703
rect 20680 36672 23581 36700
rect 20680 36660 20686 36672
rect 23569 36669 23581 36672
rect 23615 36669 23627 36703
rect 36648 36700 36676 36731
rect 23569 36663 23627 36669
rect 36004 36672 36676 36700
rect 36004 36641 36032 36672
rect 14277 36635 14335 36641
rect 14277 36601 14289 36635
rect 14323 36601 14335 36635
rect 14277 36595 14335 36601
rect 35989 36635 36047 36641
rect 35989 36601 36001 36635
rect 36035 36601 36047 36635
rect 35989 36595 36047 36601
rect 2869 36567 2927 36573
rect 2869 36533 2881 36567
rect 2915 36564 2927 36567
rect 5718 36564 5724 36576
rect 2915 36536 5724 36564
rect 2915 36533 2927 36536
rect 2869 36527 2927 36533
rect 5718 36524 5724 36536
rect 5776 36524 5782 36576
rect 33134 36524 33140 36576
rect 33192 36564 33198 36576
rect 35345 36567 35403 36573
rect 35345 36564 35357 36567
rect 33192 36536 35357 36564
rect 33192 36524 33198 36536
rect 35345 36533 35357 36536
rect 35391 36533 35403 36567
rect 35345 36527 35403 36533
rect 37918 36524 37924 36576
rect 37976 36564 37982 36576
rect 38197 36567 38255 36573
rect 38197 36564 38209 36567
rect 37976 36536 38209 36564
rect 37976 36524 37982 36536
rect 38197 36533 38209 36536
rect 38243 36533 38255 36567
rect 38197 36527 38255 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1762 36360 1768 36372
rect 1723 36332 1768 36360
rect 1762 36320 1768 36332
rect 1820 36320 1826 36372
rect 9122 36320 9128 36372
rect 9180 36360 9186 36372
rect 18598 36360 18604 36372
rect 9180 36332 18604 36360
rect 9180 36320 9186 36332
rect 18598 36320 18604 36332
rect 18656 36320 18662 36372
rect 35621 36363 35679 36369
rect 35621 36329 35633 36363
rect 35667 36360 35679 36363
rect 36170 36360 36176 36372
rect 35667 36332 36176 36360
rect 35667 36329 35679 36332
rect 35621 36323 35679 36329
rect 36170 36320 36176 36332
rect 36228 36320 36234 36372
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 37240 36332 37473 36360
rect 37240 36320 37246 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 36633 36295 36691 36301
rect 36633 36261 36645 36295
rect 36679 36261 36691 36295
rect 36633 36255 36691 36261
rect 36648 36224 36676 36255
rect 36648 36196 38056 36224
rect 1578 36156 1584 36168
rect 1539 36128 1584 36156
rect 1578 36116 1584 36128
rect 1636 36116 1642 36168
rect 2501 36159 2559 36165
rect 2501 36125 2513 36159
rect 2547 36156 2559 36159
rect 2774 36156 2780 36168
rect 2547 36128 2780 36156
rect 2547 36125 2559 36128
rect 2501 36119 2559 36125
rect 2774 36116 2780 36128
rect 2832 36116 2838 36168
rect 35526 36156 35532 36168
rect 35487 36128 35532 36156
rect 35526 36116 35532 36128
rect 35584 36116 35590 36168
rect 36814 36156 36820 36168
rect 36775 36128 36820 36156
rect 36814 36116 36820 36128
rect 36872 36116 36878 36168
rect 37274 36156 37280 36168
rect 37235 36128 37280 36156
rect 37274 36116 37280 36128
rect 37332 36116 37338 36168
rect 38028 36165 38056 36196
rect 38013 36159 38071 36165
rect 38013 36125 38025 36159
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 2317 36023 2375 36029
rect 2317 35989 2329 36023
rect 2363 36020 2375 36023
rect 6822 36020 6828 36032
rect 2363 35992 6828 36020
rect 2363 35989 2375 35992
rect 2317 35983 2375 35989
rect 6822 35980 6828 35992
rect 6880 35980 6886 36032
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 18690 35776 18696 35828
rect 18748 35816 18754 35828
rect 19426 35816 19432 35828
rect 18748 35788 19432 35816
rect 18748 35776 18754 35788
rect 19426 35776 19432 35788
rect 19484 35776 19490 35828
rect 1581 35683 1639 35689
rect 1581 35649 1593 35683
rect 1627 35680 1639 35683
rect 4614 35680 4620 35692
rect 1627 35652 4620 35680
rect 1627 35649 1639 35652
rect 1581 35643 1639 35649
rect 4614 35640 4620 35652
rect 4672 35640 4678 35692
rect 37826 35640 37832 35692
rect 37884 35680 37890 35692
rect 38013 35683 38071 35689
rect 38013 35680 38025 35683
rect 37884 35652 38025 35680
rect 37884 35640 37890 35652
rect 38013 35649 38025 35652
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 1762 35476 1768 35488
rect 1723 35448 1768 35476
rect 1762 35436 1768 35448
rect 1820 35436 1826 35488
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 22278 35164 22284 35216
rect 22336 35204 22342 35216
rect 37274 35204 37280 35216
rect 22336 35176 37280 35204
rect 22336 35164 22342 35176
rect 37274 35164 37280 35176
rect 37332 35164 37338 35216
rect 1762 35068 1768 35080
rect 1723 35040 1768 35068
rect 1762 35028 1768 35040
rect 1820 35028 1826 35080
rect 37366 35028 37372 35080
rect 37424 35068 37430 35080
rect 37645 35071 37703 35077
rect 37645 35068 37657 35071
rect 37424 35040 37657 35068
rect 37424 35028 37430 35040
rect 37645 35037 37657 35040
rect 37691 35037 37703 35071
rect 37645 35031 37703 35037
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 4062 34932 4068 34944
rect 1627 34904 4068 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 4062 34892 4068 34904
rect 4120 34892 4126 34944
rect 37458 34932 37464 34944
rect 37419 34904 37464 34932
rect 37458 34892 37464 34904
rect 37516 34892 37522 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 14185 34731 14243 34737
rect 14185 34697 14197 34731
rect 14231 34728 14243 34731
rect 15378 34728 15384 34740
rect 14231 34700 15384 34728
rect 14231 34697 14243 34700
rect 14185 34691 14243 34697
rect 15378 34688 15384 34700
rect 15436 34688 15442 34740
rect 35253 34731 35311 34737
rect 35253 34697 35265 34731
rect 35299 34728 35311 34731
rect 35989 34731 36047 34737
rect 35299 34700 35894 34728
rect 35299 34697 35311 34700
rect 35253 34691 35311 34697
rect 35866 34660 35894 34700
rect 35989 34697 36001 34731
rect 36035 34728 36047 34731
rect 36814 34728 36820 34740
rect 36035 34700 36820 34728
rect 36035 34697 36047 34700
rect 35989 34691 36047 34697
rect 36814 34688 36820 34700
rect 36872 34688 36878 34740
rect 35866 34632 38056 34660
rect 13906 34552 13912 34604
rect 13964 34592 13970 34604
rect 14369 34595 14427 34601
rect 14369 34592 14381 34595
rect 13964 34564 14381 34592
rect 13964 34552 13970 34564
rect 14369 34561 14381 34564
rect 14415 34561 14427 34595
rect 35434 34592 35440 34604
rect 35395 34564 35440 34592
rect 14369 34555 14427 34561
rect 35434 34552 35440 34564
rect 35492 34552 35498 34604
rect 35897 34595 35955 34601
rect 35897 34561 35909 34595
rect 35943 34592 35955 34595
rect 35986 34592 35992 34604
rect 35943 34564 35992 34592
rect 35943 34561 35955 34564
rect 35897 34555 35955 34561
rect 35986 34552 35992 34564
rect 36044 34552 36050 34604
rect 38028 34601 38056 34632
rect 38013 34595 38071 34601
rect 38013 34561 38025 34595
rect 38059 34561 38071 34595
rect 38013 34555 38071 34561
rect 21358 34484 21364 34536
rect 21416 34524 21422 34536
rect 24578 34524 24584 34536
rect 21416 34496 24584 34524
rect 21416 34484 21422 34496
rect 24578 34484 24584 34496
rect 24636 34484 24642 34536
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 18969 33643 19027 33649
rect 18969 33640 18981 33643
rect 6886 33612 18981 33640
rect 1581 33507 1639 33513
rect 1581 33473 1593 33507
rect 1627 33504 1639 33507
rect 6886 33504 6914 33612
rect 18969 33609 18981 33612
rect 19015 33609 19027 33643
rect 18969 33603 19027 33609
rect 19150 33504 19156 33516
rect 1627 33476 6914 33504
rect 19111 33476 19156 33504
rect 1627 33473 1639 33476
rect 1581 33467 1639 33473
rect 19150 33464 19156 33476
rect 19208 33464 19214 33516
rect 1762 33368 1768 33380
rect 1723 33340 1768 33368
rect 1762 33328 1768 33340
rect 1820 33328 1826 33380
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 5718 32892 5724 32904
rect 5679 32864 5724 32892
rect 5718 32852 5724 32864
rect 5776 32852 5782 32904
rect 23753 32895 23811 32901
rect 23753 32861 23765 32895
rect 23799 32892 23811 32895
rect 28534 32892 28540 32904
rect 23799 32864 28540 32892
rect 23799 32861 23811 32864
rect 23753 32855 23811 32861
rect 28534 32852 28540 32864
rect 28592 32852 28598 32904
rect 36446 32852 36452 32904
rect 36504 32892 36510 32904
rect 38013 32895 38071 32901
rect 38013 32892 38025 32895
rect 36504 32864 38025 32892
rect 36504 32852 36510 32864
rect 38013 32861 38025 32864
rect 38059 32861 38071 32895
rect 38013 32855 38071 32861
rect 5813 32759 5871 32765
rect 5813 32725 5825 32759
rect 5859 32756 5871 32759
rect 6638 32756 6644 32768
rect 5859 32728 6644 32756
rect 5859 32725 5871 32728
rect 5813 32719 5871 32725
rect 6638 32716 6644 32728
rect 6696 32716 6702 32768
rect 17770 32716 17776 32768
rect 17828 32756 17834 32768
rect 23845 32759 23903 32765
rect 23845 32756 23857 32759
rect 17828 32728 23857 32756
rect 17828 32716 17834 32728
rect 23845 32725 23857 32728
rect 23891 32725 23903 32759
rect 38194 32756 38200 32768
rect 38155 32728 38200 32756
rect 23845 32719 23903 32725
rect 38194 32716 38200 32728
rect 38252 32716 38258 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 5810 32376 5816 32428
rect 5868 32416 5874 32428
rect 9033 32419 9091 32425
rect 9033 32416 9045 32419
rect 5868 32388 9045 32416
rect 5868 32376 5874 32388
rect 9033 32385 9045 32388
rect 9079 32385 9091 32419
rect 9033 32379 9091 32385
rect 33226 32376 33232 32428
rect 33284 32416 33290 32428
rect 38013 32419 38071 32425
rect 38013 32416 38025 32419
rect 33284 32388 38025 32416
rect 33284 32376 33290 32388
rect 38013 32385 38025 32388
rect 38059 32385 38071 32419
rect 38013 32379 38071 32385
rect 1578 32348 1584 32360
rect 1539 32320 1584 32348
rect 1578 32308 1584 32320
rect 1636 32308 1642 32360
rect 1857 32351 1915 32357
rect 1857 32317 1869 32351
rect 1903 32348 1915 32351
rect 9306 32348 9312 32360
rect 1903 32320 9312 32348
rect 1903 32317 1915 32320
rect 1857 32311 1915 32317
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 9122 32212 9128 32224
rect 9083 32184 9128 32212
rect 9122 32172 9128 32184
rect 9180 32172 9186 32224
rect 38194 32212 38200 32224
rect 38155 32184 38200 32212
rect 38194 32172 38200 32184
rect 38252 32172 38258 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 4525 32011 4583 32017
rect 4525 31977 4537 32011
rect 4571 32008 4583 32011
rect 4614 32008 4620 32020
rect 4571 31980 4620 32008
rect 4571 31977 4583 31980
rect 4525 31971 4583 31977
rect 4614 31968 4620 31980
rect 4672 31968 4678 32020
rect 7469 32011 7527 32017
rect 7469 31977 7481 32011
rect 7515 32008 7527 32011
rect 7834 32008 7840 32020
rect 7515 31980 7840 32008
rect 7515 31977 7527 31980
rect 7469 31971 7527 31977
rect 7834 31968 7840 31980
rect 7892 31968 7898 32020
rect 17402 31968 17408 32020
rect 17460 32008 17466 32020
rect 24673 32011 24731 32017
rect 24673 32008 24685 32011
rect 17460 31980 24685 32008
rect 17460 31968 17466 31980
rect 24673 31977 24685 31980
rect 24719 31977 24731 32011
rect 24673 31971 24731 31977
rect 9030 31900 9036 31952
rect 9088 31940 9094 31952
rect 9217 31943 9275 31949
rect 9217 31940 9229 31943
rect 9088 31912 9229 31940
rect 9088 31900 9094 31912
rect 9217 31909 9229 31912
rect 9263 31909 9275 31943
rect 9217 31903 9275 31909
rect 20254 31900 20260 31952
rect 20312 31940 20318 31952
rect 21821 31943 21879 31949
rect 21821 31940 21833 31943
rect 20312 31912 21833 31940
rect 20312 31900 20318 31912
rect 21821 31909 21833 31912
rect 21867 31909 21879 31943
rect 21821 31903 21879 31909
rect 6546 31832 6552 31884
rect 6604 31872 6610 31884
rect 6604 31844 9168 31872
rect 6604 31832 6610 31844
rect 1581 31807 1639 31813
rect 1581 31773 1593 31807
rect 1627 31804 1639 31807
rect 4614 31804 4620 31816
rect 1627 31776 4620 31804
rect 1627 31773 1639 31776
rect 1581 31767 1639 31773
rect 4614 31764 4620 31776
rect 4672 31764 4678 31816
rect 4709 31807 4767 31813
rect 4709 31773 4721 31807
rect 4755 31804 4767 31807
rect 6730 31804 6736 31816
rect 4755 31776 6736 31804
rect 4755 31773 4767 31776
rect 4709 31767 4767 31773
rect 6730 31764 6736 31776
rect 6788 31764 6794 31816
rect 7650 31804 7656 31816
rect 7611 31776 7656 31804
rect 7650 31764 7656 31776
rect 7708 31764 7714 31816
rect 9140 31813 9168 31844
rect 14182 31832 14188 31884
rect 14240 31872 14246 31884
rect 15933 31875 15991 31881
rect 15933 31872 15945 31875
rect 14240 31844 15945 31872
rect 14240 31832 14246 31844
rect 15933 31841 15945 31844
rect 15979 31841 15991 31875
rect 25314 31872 25320 31884
rect 15933 31835 15991 31841
rect 21744 31844 25320 31872
rect 9125 31807 9183 31813
rect 9125 31773 9137 31807
rect 9171 31773 9183 31807
rect 9125 31767 9183 31773
rect 15841 31807 15899 31813
rect 15841 31773 15853 31807
rect 15887 31804 15899 31807
rect 19334 31804 19340 31816
rect 15887 31776 19340 31804
rect 15887 31773 15899 31776
rect 15841 31767 15899 31773
rect 19334 31764 19340 31776
rect 19392 31764 19398 31816
rect 21744 31813 21772 31844
rect 25314 31832 25320 31844
rect 25372 31832 25378 31884
rect 21729 31807 21787 31813
rect 21729 31773 21741 31807
rect 21775 31773 21787 31807
rect 21729 31767 21787 31773
rect 24581 31807 24639 31813
rect 24581 31773 24593 31807
rect 24627 31804 24639 31807
rect 28626 31804 28632 31816
rect 24627 31776 28632 31804
rect 24627 31773 24639 31776
rect 24581 31767 24639 31773
rect 28626 31764 28632 31776
rect 28684 31764 28690 31816
rect 1762 31668 1768 31680
rect 1723 31640 1768 31668
rect 1762 31628 1768 31640
rect 1820 31628 1826 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 7469 31467 7527 31473
rect 7469 31433 7481 31467
rect 7515 31464 7527 31467
rect 7650 31464 7656 31476
rect 7515 31436 7656 31464
rect 7515 31433 7527 31436
rect 7469 31427 7527 31433
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 7374 31328 7380 31340
rect 7335 31300 7380 31328
rect 7374 31288 7380 31300
rect 7432 31288 7438 31340
rect 23937 31331 23995 31337
rect 23937 31297 23949 31331
rect 23983 31328 23995 31331
rect 26234 31328 26240 31340
rect 23983 31300 26240 31328
rect 23983 31297 23995 31300
rect 23937 31291 23995 31297
rect 26234 31288 26240 31300
rect 26292 31288 26298 31340
rect 28629 31331 28687 31337
rect 28629 31297 28641 31331
rect 28675 31328 28687 31331
rect 37458 31328 37464 31340
rect 28675 31300 37464 31328
rect 28675 31297 28687 31300
rect 28629 31291 28687 31297
rect 37458 31288 37464 31300
rect 37516 31288 37522 31340
rect 20346 31084 20352 31136
rect 20404 31124 20410 31136
rect 24029 31127 24087 31133
rect 24029 31124 24041 31127
rect 20404 31096 24041 31124
rect 20404 31084 20410 31096
rect 24029 31093 24041 31096
rect 24075 31093 24087 31127
rect 24029 31087 24087 31093
rect 26694 31084 26700 31136
rect 26752 31124 26758 31136
rect 28721 31127 28779 31133
rect 28721 31124 28733 31127
rect 26752 31096 28733 31124
rect 26752 31084 26758 31096
rect 28721 31093 28733 31096
rect 28767 31093 28779 31127
rect 28721 31087 28779 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 4062 30676 4068 30728
rect 4120 30716 4126 30728
rect 4985 30719 5043 30725
rect 4985 30716 4997 30719
rect 4120 30688 4997 30716
rect 4120 30676 4126 30688
rect 4985 30685 4997 30688
rect 5031 30685 5043 30719
rect 9398 30716 9404 30728
rect 9359 30688 9404 30716
rect 4985 30679 5043 30685
rect 9398 30676 9404 30688
rect 9456 30676 9462 30728
rect 22097 30719 22155 30725
rect 22097 30685 22109 30719
rect 22143 30716 22155 30719
rect 27154 30716 27160 30728
rect 22143 30688 27160 30716
rect 22143 30685 22155 30688
rect 22097 30679 22155 30685
rect 27154 30676 27160 30688
rect 27212 30676 27218 30728
rect 38286 30716 38292 30728
rect 38247 30688 38292 30716
rect 38286 30676 38292 30688
rect 38344 30676 38350 30728
rect 1854 30608 1860 30660
rect 1912 30648 1918 30660
rect 20073 30651 20131 30657
rect 20073 30648 20085 30651
rect 1912 30620 20085 30648
rect 1912 30608 1918 30620
rect 20073 30617 20085 30620
rect 20119 30617 20131 30651
rect 20073 30611 20131 30617
rect 20257 30651 20315 30657
rect 20257 30617 20269 30651
rect 20303 30648 20315 30651
rect 33686 30648 33692 30660
rect 20303 30620 33692 30648
rect 20303 30617 20315 30620
rect 20257 30611 20315 30617
rect 33686 30608 33692 30620
rect 33744 30608 33750 30660
rect 5077 30583 5135 30589
rect 5077 30549 5089 30583
rect 5123 30580 5135 30583
rect 8570 30580 8576 30592
rect 5123 30552 8576 30580
rect 5123 30549 5135 30552
rect 5077 30543 5135 30549
rect 8570 30540 8576 30552
rect 8628 30540 8634 30592
rect 9493 30583 9551 30589
rect 9493 30549 9505 30583
rect 9539 30580 9551 30583
rect 11330 30580 11336 30592
rect 9539 30552 11336 30580
rect 9539 30549 9551 30552
rect 9493 30543 9551 30549
rect 11330 30540 11336 30552
rect 11388 30540 11394 30592
rect 17126 30540 17132 30592
rect 17184 30580 17190 30592
rect 22189 30583 22247 30589
rect 22189 30580 22201 30583
rect 17184 30552 22201 30580
rect 17184 30540 17190 30552
rect 22189 30549 22201 30552
rect 22235 30549 22247 30583
rect 22189 30543 22247 30549
rect 36998 30540 37004 30592
rect 37056 30580 37062 30592
rect 38105 30583 38163 30589
rect 38105 30580 38117 30583
rect 37056 30552 38117 30580
rect 37056 30540 37062 30552
rect 38105 30549 38117 30552
rect 38151 30549 38163 30583
rect 38105 30543 38163 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 33042 30308 33048 30320
rect 25884 30280 33048 30308
rect 1581 30243 1639 30249
rect 1581 30209 1593 30243
rect 1627 30240 1639 30243
rect 5442 30240 5448 30252
rect 1627 30212 5448 30240
rect 1627 30209 1639 30212
rect 1581 30203 1639 30209
rect 5442 30200 5448 30212
rect 5500 30200 5506 30252
rect 12342 30240 12348 30252
rect 12303 30212 12348 30240
rect 12342 30200 12348 30212
rect 12400 30200 12406 30252
rect 25884 30249 25912 30280
rect 33042 30268 33048 30280
rect 33100 30268 33106 30320
rect 25869 30243 25927 30249
rect 25869 30209 25881 30243
rect 25915 30209 25927 30243
rect 25869 30203 25927 30209
rect 27157 30243 27215 30249
rect 27157 30209 27169 30243
rect 27203 30240 27215 30243
rect 33134 30240 33140 30252
rect 27203 30212 33140 30240
rect 27203 30209 27215 30212
rect 27157 30203 27215 30209
rect 33134 30200 33140 30212
rect 33192 30200 33198 30252
rect 17218 30064 17224 30116
rect 17276 30104 17282 30116
rect 27249 30107 27307 30113
rect 27249 30104 27261 30107
rect 17276 30076 27261 30104
rect 17276 30064 17282 30076
rect 27249 30073 27261 30076
rect 27295 30073 27307 30107
rect 27249 30067 27307 30073
rect 1762 30036 1768 30048
rect 1723 30008 1768 30036
rect 1762 29996 1768 30008
rect 1820 29996 1826 30048
rect 12434 29996 12440 30048
rect 12492 30036 12498 30048
rect 12492 30008 12537 30036
rect 12492 29996 12498 30008
rect 18230 29996 18236 30048
rect 18288 30036 18294 30048
rect 25961 30039 26019 30045
rect 25961 30036 25973 30039
rect 18288 30008 25973 30036
rect 18288 29996 18294 30008
rect 25961 30005 25973 30008
rect 26007 30005 26019 30039
rect 25961 29999 26019 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 6730 29832 6736 29844
rect 6691 29804 6736 29832
rect 6730 29792 6736 29804
rect 6788 29792 6794 29844
rect 3970 29656 3976 29708
rect 4028 29696 4034 29708
rect 4028 29668 9168 29696
rect 4028 29656 4034 29668
rect 6641 29631 6699 29637
rect 6641 29597 6653 29631
rect 6687 29628 6699 29631
rect 8938 29628 8944 29640
rect 6687 29600 8944 29628
rect 6687 29597 6699 29600
rect 6641 29591 6699 29597
rect 8938 29588 8944 29600
rect 8996 29588 9002 29640
rect 9140 29637 9168 29668
rect 9125 29631 9183 29637
rect 9125 29597 9137 29631
rect 9171 29597 9183 29631
rect 9125 29591 9183 29597
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 35894 29628 35900 29640
rect 20036 29600 35900 29628
rect 20036 29588 20042 29600
rect 35894 29588 35900 29600
rect 35952 29588 35958 29640
rect 38102 29560 38108 29572
rect 38063 29532 38108 29560
rect 38102 29520 38108 29532
rect 38160 29520 38166 29572
rect 9217 29495 9275 29501
rect 9217 29461 9229 29495
rect 9263 29492 9275 29495
rect 10594 29492 10600 29504
rect 9263 29464 10600 29492
rect 9263 29461 9275 29464
rect 9217 29455 9275 29461
rect 10594 29452 10600 29464
rect 10652 29452 10658 29504
rect 37734 29452 37740 29504
rect 37792 29492 37798 29504
rect 38197 29495 38255 29501
rect 38197 29492 38209 29495
rect 37792 29464 38209 29492
rect 37792 29452 37798 29464
rect 38197 29461 38209 29464
rect 38243 29461 38255 29495
rect 38197 29455 38255 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 4433 29291 4491 29297
rect 4433 29257 4445 29291
rect 4479 29288 4491 29291
rect 4614 29288 4620 29300
rect 4479 29260 4620 29288
rect 4479 29257 4491 29260
rect 4433 29251 4491 29257
rect 4614 29248 4620 29260
rect 4672 29248 4678 29300
rect 33226 29288 33232 29300
rect 33187 29260 33232 29288
rect 33226 29248 33232 29260
rect 33284 29248 33290 29300
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 4617 29155 4675 29161
rect 4617 29121 4629 29155
rect 4663 29152 4675 29155
rect 5902 29152 5908 29164
rect 4663 29124 5908 29152
rect 4663 29121 4675 29124
rect 4617 29115 4675 29121
rect 5902 29112 5908 29124
rect 5960 29112 5966 29164
rect 6822 29112 6828 29164
rect 6880 29152 6886 29164
rect 7101 29155 7159 29161
rect 7101 29152 7113 29155
rect 6880 29124 7113 29152
rect 6880 29112 6886 29124
rect 7101 29121 7113 29124
rect 7147 29121 7159 29155
rect 7101 29115 7159 29121
rect 31754 29112 31760 29164
rect 31812 29152 31818 29164
rect 33413 29155 33471 29161
rect 33413 29152 33425 29155
rect 31812 29124 33425 29152
rect 31812 29112 31818 29124
rect 33413 29121 33425 29124
rect 33459 29121 33471 29155
rect 33413 29115 33471 29121
rect 1581 29019 1639 29025
rect 1581 28985 1593 29019
rect 1627 29016 1639 29019
rect 2682 29016 2688 29028
rect 1627 28988 2688 29016
rect 1627 28985 1639 28988
rect 1581 28979 1639 28985
rect 2682 28976 2688 28988
rect 2740 28976 2746 29028
rect 6822 28976 6828 29028
rect 6880 29016 6886 29028
rect 7193 29019 7251 29025
rect 7193 29016 7205 29019
rect 6880 28988 7205 29016
rect 6880 28976 6886 28988
rect 7193 28985 7205 28988
rect 7239 28985 7251 29019
rect 7193 28979 7251 28985
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 15105 28543 15163 28549
rect 15105 28509 15117 28543
rect 15151 28540 15163 28543
rect 15562 28540 15568 28552
rect 15151 28512 15568 28540
rect 15151 28509 15163 28512
rect 15105 28503 15163 28509
rect 15562 28500 15568 28512
rect 15620 28500 15626 28552
rect 26237 28543 26295 28549
rect 26237 28509 26249 28543
rect 26283 28540 26295 28543
rect 35434 28540 35440 28552
rect 26283 28512 35440 28540
rect 26283 28509 26295 28512
rect 26237 28503 26295 28509
rect 35434 28500 35440 28512
rect 35492 28500 35498 28552
rect 2866 28432 2872 28484
rect 2924 28472 2930 28484
rect 20714 28472 20720 28484
rect 2924 28444 20720 28472
rect 2924 28432 2930 28444
rect 20714 28432 20720 28444
rect 20772 28432 20778 28484
rect 15197 28407 15255 28413
rect 15197 28373 15209 28407
rect 15243 28404 15255 28407
rect 15746 28404 15752 28416
rect 15243 28376 15752 28404
rect 15243 28373 15255 28376
rect 15197 28367 15255 28373
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 24854 28364 24860 28416
rect 24912 28404 24918 28416
rect 26329 28407 26387 28413
rect 26329 28404 26341 28407
rect 24912 28376 26341 28404
rect 24912 28364 24918 28376
rect 26329 28373 26341 28376
rect 26375 28373 26387 28407
rect 26329 28367 26387 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 32309 28203 32367 28209
rect 32309 28169 32321 28203
rect 32355 28200 32367 28203
rect 36446 28200 36452 28212
rect 32355 28172 36452 28200
rect 32355 28169 32367 28172
rect 32309 28163 32367 28169
rect 36446 28160 36452 28172
rect 36504 28160 36510 28212
rect 15194 28092 15200 28144
rect 15252 28132 15258 28144
rect 17037 28135 17095 28141
rect 17037 28132 17049 28135
rect 15252 28104 17049 28132
rect 15252 28092 15258 28104
rect 17037 28101 17049 28104
rect 17083 28101 17095 28135
rect 17037 28095 17095 28101
rect 1394 28024 1400 28076
rect 1452 28064 1458 28076
rect 1765 28067 1823 28073
rect 1765 28064 1777 28067
rect 1452 28036 1777 28064
rect 1452 28024 1458 28036
rect 1765 28033 1777 28036
rect 1811 28033 1823 28067
rect 1765 28027 1823 28033
rect 18417 28067 18475 28073
rect 18417 28033 18429 28067
rect 18463 28064 18475 28067
rect 19150 28064 19156 28076
rect 18463 28036 19156 28064
rect 18463 28033 18475 28036
rect 18417 28027 18475 28033
rect 19150 28024 19156 28036
rect 19208 28024 19214 28076
rect 24026 28024 24032 28076
rect 24084 28064 24090 28076
rect 29273 28067 29331 28073
rect 29273 28064 29285 28067
rect 24084 28036 29285 28064
rect 24084 28024 24090 28036
rect 29273 28033 29285 28036
rect 29319 28033 29331 28067
rect 29273 28027 29331 28033
rect 29365 28067 29423 28073
rect 29365 28033 29377 28067
rect 29411 28064 29423 28067
rect 32493 28067 32551 28073
rect 32493 28064 32505 28067
rect 29411 28036 32505 28064
rect 29411 28033 29423 28036
rect 29365 28027 29423 28033
rect 32493 28033 32505 28036
rect 32539 28033 32551 28067
rect 38286 28064 38292 28076
rect 38247 28036 38292 28064
rect 32493 28027 32551 28033
rect 38286 28024 38292 28036
rect 38344 28024 38350 28076
rect 16945 27999 17003 28005
rect 16945 27965 16957 27999
rect 16991 27996 17003 27999
rect 16991 27968 18184 27996
rect 16991 27965 17003 27968
rect 16945 27959 17003 27965
rect 17497 27931 17555 27937
rect 17497 27897 17509 27931
rect 17543 27928 17555 27931
rect 17954 27928 17960 27940
rect 17543 27900 17960 27928
rect 17543 27897 17555 27900
rect 17497 27891 17555 27897
rect 17954 27888 17960 27900
rect 18012 27888 18018 27940
rect 18156 27872 18184 27968
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 5166 27860 5172 27872
rect 1627 27832 5172 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 5166 27820 5172 27832
rect 5224 27820 5230 27872
rect 11238 27820 11244 27872
rect 11296 27860 11302 27872
rect 14182 27860 14188 27872
rect 11296 27832 14188 27860
rect 11296 27820 11302 27832
rect 14182 27820 14188 27832
rect 14240 27820 14246 27872
rect 18138 27820 18144 27872
rect 18196 27860 18202 27872
rect 18509 27863 18567 27869
rect 18509 27860 18521 27863
rect 18196 27832 18521 27860
rect 18196 27820 18202 27832
rect 18509 27829 18521 27832
rect 18555 27829 18567 27863
rect 18509 27823 18567 27829
rect 36078 27820 36084 27872
rect 36136 27860 36142 27872
rect 38105 27863 38163 27869
rect 38105 27860 38117 27863
rect 36136 27832 38117 27860
rect 36136 27820 36142 27832
rect 38105 27829 38117 27832
rect 38151 27829 38163 27863
rect 38105 27823 38163 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 28445 27591 28503 27597
rect 28445 27557 28457 27591
rect 28491 27588 28503 27591
rect 31754 27588 31760 27600
rect 28491 27560 31760 27588
rect 28491 27557 28503 27560
rect 28445 27551 28503 27557
rect 31754 27548 31760 27560
rect 31812 27548 31818 27600
rect 5994 27480 6000 27532
rect 6052 27520 6058 27532
rect 12342 27520 12348 27532
rect 6052 27492 12348 27520
rect 6052 27480 6058 27492
rect 12342 27480 12348 27492
rect 12400 27520 12406 27532
rect 12400 27492 12480 27520
rect 12400 27480 12406 27492
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27421 1639 27455
rect 1581 27415 1639 27421
rect 2317 27455 2375 27461
rect 2317 27421 2329 27455
rect 2363 27452 2375 27455
rect 2406 27452 2412 27464
rect 2363 27424 2412 27452
rect 2363 27421 2375 27424
rect 2317 27415 2375 27421
rect 1596 27384 1624 27415
rect 2406 27412 2412 27424
rect 2464 27412 2470 27464
rect 11609 27455 11667 27461
rect 11609 27421 11621 27455
rect 11655 27452 11667 27455
rect 11974 27452 11980 27464
rect 11655 27424 11980 27452
rect 11655 27421 11667 27424
rect 11609 27415 11667 27421
rect 11974 27412 11980 27424
rect 12032 27412 12038 27464
rect 12452 27461 12480 27492
rect 12912 27492 13676 27520
rect 12912 27461 12940 27492
rect 13648 27464 13676 27492
rect 12437 27455 12495 27461
rect 12437 27421 12449 27455
rect 12483 27421 12495 27455
rect 12437 27415 12495 27421
rect 12897 27455 12955 27461
rect 12897 27421 12909 27455
rect 12943 27421 12955 27455
rect 13538 27452 13544 27464
rect 13499 27424 13544 27452
rect 12897 27415 12955 27421
rect 13538 27412 13544 27424
rect 13596 27412 13602 27464
rect 13630 27412 13636 27464
rect 13688 27452 13694 27464
rect 14277 27455 14335 27461
rect 14277 27452 14289 27455
rect 13688 27424 14289 27452
rect 13688 27412 13694 27424
rect 14277 27421 14289 27424
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 26234 27412 26240 27464
rect 26292 27452 26298 27464
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 26292 27424 28365 27452
rect 26292 27412 26298 27424
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 28353 27415 28411 27421
rect 35894 27412 35900 27464
rect 35952 27452 35958 27464
rect 38013 27455 38071 27461
rect 38013 27452 38025 27455
rect 35952 27424 38025 27452
rect 35952 27412 35958 27424
rect 38013 27421 38025 27424
rect 38059 27421 38071 27455
rect 38013 27415 38071 27421
rect 5258 27384 5264 27396
rect 1596 27356 5264 27384
rect 5258 27344 5264 27356
rect 5316 27344 5322 27396
rect 9766 27344 9772 27396
rect 9824 27384 9830 27396
rect 14458 27384 14464 27396
rect 9824 27356 14464 27384
rect 9824 27344 9830 27356
rect 14458 27344 14464 27356
rect 14516 27344 14522 27396
rect 1762 27316 1768 27328
rect 1723 27288 1768 27316
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 2409 27319 2467 27325
rect 2409 27285 2421 27319
rect 2455 27316 2467 27319
rect 2498 27316 2504 27328
rect 2455 27288 2504 27316
rect 2455 27285 2467 27288
rect 2409 27279 2467 27285
rect 2498 27276 2504 27288
rect 2556 27276 2562 27328
rect 11054 27276 11060 27328
rect 11112 27316 11118 27328
rect 11425 27319 11483 27325
rect 11425 27316 11437 27319
rect 11112 27288 11437 27316
rect 11112 27276 11118 27288
rect 11425 27285 11437 27288
rect 11471 27285 11483 27319
rect 12250 27316 12256 27328
rect 12211 27288 12256 27316
rect 11425 27279 11483 27285
rect 12250 27276 12256 27288
rect 12308 27276 12314 27328
rect 12618 27276 12624 27328
rect 12676 27316 12682 27328
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 12676 27288 13001 27316
rect 12676 27276 12682 27288
rect 12989 27285 13001 27288
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13446 27276 13452 27328
rect 13504 27316 13510 27328
rect 13633 27319 13691 27325
rect 13633 27316 13645 27319
rect 13504 27288 13645 27316
rect 13504 27276 13510 27288
rect 13633 27285 13645 27288
rect 13679 27285 13691 27319
rect 14366 27316 14372 27328
rect 14327 27288 14372 27316
rect 13633 27279 13691 27285
rect 14366 27276 14372 27288
rect 14424 27276 14430 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 5902 27112 5908 27124
rect 5863 27084 5908 27112
rect 5902 27072 5908 27084
rect 5960 27072 5966 27124
rect 8202 27072 8208 27124
rect 8260 27112 8266 27124
rect 14553 27115 14611 27121
rect 8260 27084 11744 27112
rect 8260 27072 8266 27084
rect 6825 27047 6883 27053
rect 6825 27013 6837 27047
rect 6871 27044 6883 27047
rect 8757 27047 8815 27053
rect 8757 27044 8769 27047
rect 6871 27016 8769 27044
rect 6871 27013 6883 27016
rect 6825 27007 6883 27013
rect 8757 27013 8769 27016
rect 8803 27013 8815 27047
rect 8757 27007 8815 27013
rect 8938 27004 8944 27056
rect 8996 27044 9002 27056
rect 9309 27047 9367 27053
rect 9309 27044 9321 27047
rect 8996 27016 9321 27044
rect 8996 27004 9002 27016
rect 9309 27013 9321 27016
rect 9355 27013 9367 27047
rect 9309 27007 9367 27013
rect 1854 26976 1860 26988
rect 1815 26948 1860 26976
rect 1854 26936 1860 26948
rect 1912 26936 1918 26988
rect 2314 26936 2320 26988
rect 2372 26976 2378 26988
rect 2501 26979 2559 26985
rect 2501 26976 2513 26979
rect 2372 26948 2513 26976
rect 2372 26936 2378 26948
rect 2501 26945 2513 26948
rect 2547 26945 2559 26979
rect 2501 26939 2559 26945
rect 3145 26979 3203 26985
rect 3145 26945 3157 26979
rect 3191 26945 3203 26979
rect 5810 26976 5816 26988
rect 5771 26948 5816 26976
rect 3145 26939 3203 26945
rect 2516 26840 2544 26939
rect 3160 26908 3188 26939
rect 5810 26936 5816 26948
rect 5868 26936 5874 26988
rect 6454 26936 6460 26988
rect 6512 26976 6518 26988
rect 6733 26979 6791 26985
rect 6733 26976 6745 26979
rect 6512 26948 6745 26976
rect 6512 26936 6518 26948
rect 6733 26945 6745 26948
rect 6779 26945 6791 26979
rect 6733 26939 6791 26945
rect 7929 26979 7987 26985
rect 7929 26945 7941 26979
rect 7975 26945 7987 26979
rect 11054 26976 11060 26988
rect 11015 26948 11060 26976
rect 7929 26939 7987 26945
rect 7834 26908 7840 26920
rect 3160 26880 7840 26908
rect 7834 26868 7840 26880
rect 7892 26868 7898 26920
rect 6730 26840 6736 26852
rect 2516 26812 6736 26840
rect 6730 26800 6736 26812
rect 6788 26800 6794 26852
rect 7944 26840 7972 26939
rect 11054 26936 11060 26948
rect 11112 26936 11118 26988
rect 11716 26985 11744 27084
rect 14553 27081 14565 27115
rect 14599 27112 14611 27115
rect 15194 27112 15200 27124
rect 14599 27084 15200 27112
rect 14599 27081 14611 27084
rect 14553 27075 14611 27081
rect 15194 27072 15200 27084
rect 15252 27072 15258 27124
rect 13449 27047 13507 27053
rect 13449 27013 13461 27047
rect 13495 27044 13507 27047
rect 14366 27044 14372 27056
rect 13495 27016 14372 27044
rect 13495 27013 13507 27016
rect 13449 27007 13507 27013
rect 14366 27004 14372 27016
rect 14424 27004 14430 27056
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26945 11759 26979
rect 12342 26976 12348 26988
rect 12303 26948 12348 26976
rect 11701 26939 11759 26945
rect 12342 26936 12348 26948
rect 12400 26936 12406 26988
rect 14458 26976 14464 26988
rect 14419 26948 14464 26976
rect 14458 26936 14464 26948
rect 14516 26936 14522 26988
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26976 32367 26979
rect 36998 26976 37004 26988
rect 32355 26948 37004 26976
rect 32355 26945 32367 26948
rect 32309 26939 32367 26945
rect 36998 26936 37004 26948
rect 37056 26936 37062 26988
rect 8665 26911 8723 26917
rect 8665 26877 8677 26911
rect 8711 26908 8723 26911
rect 10870 26908 10876 26920
rect 8711 26880 10876 26908
rect 8711 26877 8723 26880
rect 8665 26871 8723 26877
rect 10870 26868 10876 26880
rect 10928 26868 10934 26920
rect 10962 26868 10968 26920
rect 11020 26908 11026 26920
rect 13357 26911 13415 26917
rect 13357 26908 13369 26911
rect 11020 26880 13369 26908
rect 11020 26868 11026 26880
rect 13357 26877 13369 26880
rect 13403 26908 13415 26911
rect 13998 26908 14004 26920
rect 13403 26880 14004 26908
rect 13403 26877 13415 26880
rect 13357 26871 13415 26877
rect 13998 26868 14004 26880
rect 14056 26868 14062 26920
rect 11793 26843 11851 26849
rect 7944 26812 11008 26840
rect 1670 26732 1676 26784
rect 1728 26772 1734 26784
rect 1949 26775 2007 26781
rect 1949 26772 1961 26775
rect 1728 26744 1961 26772
rect 1728 26732 1734 26744
rect 1949 26741 1961 26744
rect 1995 26741 2007 26775
rect 2590 26772 2596 26784
rect 2551 26744 2596 26772
rect 1949 26735 2007 26741
rect 2590 26732 2596 26744
rect 2648 26732 2654 26784
rect 3234 26772 3240 26784
rect 3195 26744 3240 26772
rect 3234 26732 3240 26744
rect 3292 26732 3298 26784
rect 8018 26772 8024 26784
rect 7979 26744 8024 26772
rect 8018 26732 8024 26744
rect 8076 26732 8082 26784
rect 10042 26732 10048 26784
rect 10100 26772 10106 26784
rect 10873 26775 10931 26781
rect 10873 26772 10885 26775
rect 10100 26744 10885 26772
rect 10100 26732 10106 26744
rect 10873 26741 10885 26744
rect 10919 26741 10931 26775
rect 10980 26772 11008 26812
rect 11793 26809 11805 26843
rect 11839 26840 11851 26843
rect 13814 26840 13820 26852
rect 11839 26812 13820 26840
rect 11839 26809 11851 26812
rect 11793 26803 11851 26809
rect 13814 26800 13820 26812
rect 13872 26800 13878 26852
rect 13906 26800 13912 26852
rect 13964 26840 13970 26852
rect 13964 26812 14009 26840
rect 13964 26800 13970 26812
rect 11974 26772 11980 26784
rect 10980 26744 11980 26772
rect 10873 26735 10931 26741
rect 11974 26732 11980 26744
rect 12032 26732 12038 26784
rect 12437 26775 12495 26781
rect 12437 26741 12449 26775
rect 12483 26772 12495 26775
rect 12526 26772 12532 26784
rect 12483 26744 12532 26772
rect 12483 26741 12495 26744
rect 12437 26735 12495 26741
rect 12526 26732 12532 26744
rect 12584 26732 12590 26784
rect 32398 26772 32404 26784
rect 32359 26744 32404 26772
rect 32398 26732 32404 26744
rect 32456 26732 32462 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 18046 26568 18052 26580
rect 9876 26540 15240 26568
rect 18007 26540 18052 26568
rect 3973 26503 4031 26509
rect 3973 26469 3985 26503
rect 4019 26500 4031 26503
rect 4062 26500 4068 26512
rect 4019 26472 4068 26500
rect 4019 26469 4031 26472
rect 3973 26463 4031 26469
rect 4062 26460 4068 26472
rect 4120 26460 4126 26512
rect 6273 26503 6331 26509
rect 6273 26469 6285 26503
rect 6319 26469 6331 26503
rect 6273 26463 6331 26469
rect 6917 26503 6975 26509
rect 6917 26469 6929 26503
rect 6963 26500 6975 26503
rect 9306 26500 9312 26512
rect 6963 26472 9312 26500
rect 6963 26469 6975 26472
rect 6917 26463 6975 26469
rect 6288 26432 6316 26463
rect 9306 26460 9312 26472
rect 9364 26460 9370 26512
rect 9876 26441 9904 26540
rect 10134 26460 10140 26512
rect 10192 26500 10198 26512
rect 10229 26503 10287 26509
rect 10229 26500 10241 26503
rect 10192 26472 10241 26500
rect 10192 26460 10198 26472
rect 10229 26469 10241 26472
rect 10275 26469 10287 26503
rect 10229 26463 10287 26469
rect 10870 26460 10876 26512
rect 10928 26500 10934 26512
rect 11333 26503 11391 26509
rect 11333 26500 11345 26503
rect 10928 26472 11345 26500
rect 10928 26460 10934 26472
rect 11333 26469 11345 26472
rect 11379 26500 11391 26503
rect 11882 26500 11888 26512
rect 11379 26472 11888 26500
rect 11379 26469 11391 26472
rect 11333 26463 11391 26469
rect 11882 26460 11888 26472
rect 11940 26460 11946 26512
rect 9861 26435 9919 26441
rect 6288 26404 7144 26432
rect 2041 26367 2099 26373
rect 2041 26333 2053 26367
rect 2087 26364 2099 26367
rect 2222 26364 2228 26376
rect 2087 26336 2228 26364
rect 2087 26333 2099 26336
rect 2041 26327 2099 26333
rect 2222 26324 2228 26336
rect 2280 26324 2286 26376
rect 2682 26364 2688 26376
rect 2643 26336 2688 26364
rect 2682 26324 2688 26336
rect 2740 26324 2746 26376
rect 4157 26367 4215 26373
rect 4157 26333 4169 26367
rect 4203 26364 4215 26367
rect 4798 26364 4804 26376
rect 4203 26336 4804 26364
rect 4203 26333 4215 26336
rect 4157 26327 4215 26333
rect 4798 26324 4804 26336
rect 4856 26324 4862 26376
rect 6454 26364 6460 26376
rect 6415 26336 6460 26364
rect 6454 26324 6460 26336
rect 6512 26324 6518 26376
rect 7116 26373 7144 26404
rect 9861 26401 9873 26435
rect 9907 26401 9919 26435
rect 10042 26432 10048 26444
rect 10003 26404 10048 26432
rect 9861 26395 9919 26401
rect 10042 26392 10048 26404
rect 10100 26392 10106 26444
rect 10962 26432 10968 26444
rect 10923 26404 10968 26432
rect 10962 26392 10968 26404
rect 11020 26392 11026 26444
rect 13906 26392 13912 26444
rect 13964 26432 13970 26444
rect 14369 26435 14427 26441
rect 14369 26432 14381 26435
rect 13964 26404 14381 26432
rect 13964 26392 13970 26404
rect 14369 26401 14381 26404
rect 14415 26401 14427 26435
rect 14369 26395 14427 26401
rect 7101 26367 7159 26373
rect 7101 26333 7113 26367
rect 7147 26333 7159 26367
rect 11146 26364 11152 26376
rect 11107 26336 11152 26364
rect 7101 26327 7159 26333
rect 11146 26324 11152 26336
rect 11204 26324 11210 26376
rect 12250 26364 12256 26376
rect 12211 26336 12256 26364
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 15212 26364 15240 26540
rect 18046 26528 18052 26540
rect 18104 26528 18110 26580
rect 35986 26568 35992 26580
rect 22066 26540 35992 26568
rect 19058 26500 19064 26512
rect 15396 26472 19064 26500
rect 15396 26441 15424 26472
rect 19058 26460 19064 26472
rect 19116 26500 19122 26512
rect 22066 26500 22094 26540
rect 35986 26528 35992 26540
rect 36044 26528 36050 26580
rect 19116 26472 22094 26500
rect 19116 26460 19122 26472
rect 34606 26460 34612 26512
rect 34664 26500 34670 26512
rect 38105 26503 38163 26509
rect 38105 26500 38117 26503
rect 34664 26472 38117 26500
rect 34664 26460 34670 26472
rect 38105 26469 38117 26472
rect 38151 26469 38163 26503
rect 38105 26463 38163 26469
rect 15381 26435 15439 26441
rect 15381 26401 15393 26435
rect 15427 26401 15439 26435
rect 16025 26435 16083 26441
rect 16025 26432 16037 26435
rect 15381 26395 15439 26401
rect 15488 26404 16037 26432
rect 15488 26364 15516 26404
rect 16025 26401 16037 26404
rect 16071 26432 16083 26435
rect 24854 26432 24860 26444
rect 16071 26404 24860 26432
rect 16071 26401 16083 26404
rect 16025 26395 16083 26401
rect 24854 26392 24860 26404
rect 24912 26392 24918 26444
rect 15212 26336 15516 26364
rect 17586 26324 17592 26376
rect 17644 26364 17650 26376
rect 18233 26367 18291 26373
rect 18233 26364 18245 26367
rect 17644 26336 18245 26364
rect 17644 26324 17650 26336
rect 18233 26333 18245 26336
rect 18279 26333 18291 26367
rect 18233 26327 18291 26333
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19613 26367 19671 26373
rect 19613 26364 19625 26367
rect 19392 26336 19625 26364
rect 19392 26324 19398 26336
rect 19613 26333 19625 26336
rect 19659 26364 19671 26367
rect 20809 26367 20867 26373
rect 20809 26364 20821 26367
rect 19659 26336 20821 26364
rect 19659 26333 19671 26336
rect 19613 26327 19671 26333
rect 20809 26333 20821 26336
rect 20855 26364 20867 26367
rect 22373 26367 22431 26373
rect 22373 26364 22385 26367
rect 20855 26336 22385 26364
rect 20855 26333 20867 26336
rect 20809 26327 20867 26333
rect 22373 26333 22385 26336
rect 22419 26333 22431 26367
rect 22373 26327 22431 26333
rect 23017 26367 23075 26373
rect 23017 26333 23029 26367
rect 23063 26333 23075 26367
rect 38286 26364 38292 26376
rect 38247 26336 38292 26364
rect 23017 26327 23075 26333
rect 2133 26299 2191 26305
rect 2133 26265 2145 26299
rect 2179 26296 2191 26299
rect 2314 26296 2320 26308
rect 2179 26268 2320 26296
rect 2179 26265 2191 26268
rect 2133 26259 2191 26265
rect 2314 26256 2320 26268
rect 2372 26256 2378 26308
rect 2777 26299 2835 26305
rect 2777 26265 2789 26299
rect 2823 26296 2835 26299
rect 2958 26296 2964 26308
rect 2823 26268 2964 26296
rect 2823 26265 2835 26268
rect 2777 26259 2835 26265
rect 2958 26256 2964 26268
rect 3016 26256 3022 26308
rect 9582 26256 9588 26308
rect 9640 26296 9646 26308
rect 14461 26299 14519 26305
rect 9640 26268 14320 26296
rect 9640 26256 9646 26268
rect 11146 26188 11152 26240
rect 11204 26228 11210 26240
rect 12069 26231 12127 26237
rect 12069 26228 12081 26231
rect 11204 26200 12081 26228
rect 11204 26188 11210 26200
rect 12069 26197 12081 26200
rect 12115 26197 12127 26231
rect 14292 26228 14320 26268
rect 14461 26265 14473 26299
rect 14507 26265 14519 26299
rect 14461 26259 14519 26265
rect 16117 26299 16175 26305
rect 16117 26265 16129 26299
rect 16163 26296 16175 26299
rect 16390 26296 16396 26308
rect 16163 26268 16396 26296
rect 16163 26265 16175 26268
rect 16117 26259 16175 26265
rect 14476 26228 14504 26259
rect 16390 26256 16396 26268
rect 16448 26256 16454 26308
rect 17037 26299 17095 26305
rect 17037 26265 17049 26299
rect 17083 26296 17095 26299
rect 17310 26296 17316 26308
rect 17083 26268 17316 26296
rect 17083 26265 17095 26268
rect 17037 26259 17095 26265
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 20162 26256 20168 26308
rect 20220 26296 20226 26308
rect 20901 26299 20959 26305
rect 20901 26296 20913 26299
rect 20220 26268 20913 26296
rect 20220 26256 20226 26268
rect 20901 26265 20913 26268
rect 20947 26265 20959 26299
rect 23032 26296 23060 26327
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 20901 26259 20959 26265
rect 22204 26268 23060 26296
rect 19426 26228 19432 26240
rect 14292 26200 14504 26228
rect 19387 26200 19432 26228
rect 12069 26191 12127 26197
rect 19426 26188 19432 26200
rect 19484 26188 19490 26240
rect 22204 26237 22232 26268
rect 22189 26231 22247 26237
rect 22189 26197 22201 26231
rect 22235 26197 22247 26231
rect 22830 26228 22836 26240
rect 22791 26200 22836 26228
rect 22189 26191 22247 26197
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 9272 25996 12572 26024
rect 9272 25984 9278 25996
rect 9493 25959 9551 25965
rect 9493 25956 9505 25959
rect 7852 25928 9505 25956
rect 1118 25848 1124 25900
rect 1176 25888 1182 25900
rect 2133 25891 2191 25897
rect 2133 25888 2145 25891
rect 1176 25860 2145 25888
rect 1176 25848 1182 25860
rect 2133 25857 2145 25860
rect 2179 25857 2191 25891
rect 3421 25891 3479 25897
rect 3421 25888 3433 25891
rect 2133 25851 2191 25857
rect 2240 25860 3433 25888
rect 1210 25780 1216 25832
rect 1268 25820 1274 25832
rect 2240 25820 2268 25860
rect 3421 25857 3433 25860
rect 3467 25857 3479 25891
rect 3421 25851 3479 25857
rect 4065 25891 4123 25897
rect 4065 25857 4077 25891
rect 4111 25857 4123 25891
rect 4890 25888 4896 25900
rect 4851 25860 4896 25888
rect 4065 25851 4123 25857
rect 1268 25792 2268 25820
rect 2777 25823 2835 25829
rect 1268 25780 1274 25792
rect 2777 25789 2789 25823
rect 2823 25820 2835 25823
rect 2866 25820 2872 25832
rect 2823 25792 2872 25820
rect 2823 25789 2835 25792
rect 2777 25783 2835 25789
rect 2866 25780 2872 25792
rect 2924 25780 2930 25832
rect 4080 25820 4108 25851
rect 4890 25848 4896 25860
rect 4948 25848 4954 25900
rect 7006 25820 7012 25832
rect 4080 25792 7012 25820
rect 7006 25780 7012 25792
rect 7064 25780 7070 25832
rect 7190 25780 7196 25832
rect 7248 25820 7254 25832
rect 7852 25829 7880 25928
rect 9493 25925 9505 25928
rect 9539 25925 9551 25959
rect 12544 25956 12572 25996
rect 13998 25984 14004 26036
rect 14056 26024 14062 26036
rect 16945 26027 17003 26033
rect 16945 26024 16957 26027
rect 14056 25996 16957 26024
rect 14056 25984 14062 25996
rect 16945 25993 16957 25996
rect 16991 25993 17003 26027
rect 16945 25987 17003 25993
rect 18598 25984 18604 26036
rect 18656 26024 18662 26036
rect 20438 26024 20444 26036
rect 18656 25996 20444 26024
rect 18656 25984 18662 25996
rect 20438 25984 20444 25996
rect 20496 25984 20502 26036
rect 18693 25959 18751 25965
rect 18693 25956 18705 25959
rect 12544 25928 14136 25956
rect 9493 25919 9551 25925
rect 8018 25888 8024 25900
rect 7979 25860 8024 25888
rect 8018 25848 8024 25860
rect 8076 25848 8082 25900
rect 9398 25888 9404 25900
rect 9359 25860 9404 25888
rect 9398 25848 9404 25860
rect 9456 25848 9462 25900
rect 10778 25888 10784 25900
rect 10739 25860 10784 25888
rect 10778 25848 10784 25860
rect 10836 25848 10842 25900
rect 12445 25889 12503 25895
rect 12445 25855 12457 25889
rect 12491 25886 12503 25889
rect 12894 25888 12900 25900
rect 12544 25886 12900 25888
rect 12491 25860 12900 25886
rect 12491 25858 12572 25860
rect 12491 25855 12503 25858
rect 12445 25849 12503 25855
rect 12894 25848 12900 25860
rect 12952 25848 12958 25900
rect 14108 25897 14136 25928
rect 16868 25928 18705 25956
rect 16868 25897 16896 25928
rect 18693 25925 18705 25928
rect 18739 25956 18751 25959
rect 18782 25956 18788 25968
rect 18739 25928 18788 25956
rect 18739 25925 18751 25928
rect 18693 25919 18751 25925
rect 18782 25916 18788 25928
rect 18840 25916 18846 25968
rect 14093 25891 14151 25897
rect 14093 25857 14105 25891
rect 14139 25857 14151 25891
rect 14093 25851 14151 25857
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25857 16911 25891
rect 16853 25851 16911 25857
rect 17957 25891 18015 25897
rect 17957 25857 17969 25891
rect 18003 25857 18015 25891
rect 17957 25851 18015 25857
rect 7837 25823 7895 25829
rect 7837 25820 7849 25823
rect 7248 25792 7849 25820
rect 7248 25780 7254 25792
rect 7837 25789 7849 25792
rect 7883 25789 7895 25823
rect 7837 25783 7895 25789
rect 7926 25780 7932 25832
rect 7984 25820 7990 25832
rect 17972 25820 18000 25851
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19521 25891 19579 25897
rect 19521 25888 19533 25891
rect 19484 25860 19533 25888
rect 19484 25848 19490 25860
rect 19521 25857 19533 25860
rect 19567 25857 19579 25891
rect 19521 25851 19579 25857
rect 19242 25820 19248 25832
rect 7984 25792 19248 25820
rect 7984 25780 7990 25792
rect 19242 25780 19248 25792
rect 19300 25780 19306 25832
rect 6730 25712 6736 25764
rect 6788 25752 6794 25764
rect 15930 25752 15936 25764
rect 6788 25724 15936 25752
rect 6788 25712 6794 25724
rect 15930 25712 15936 25724
rect 15988 25712 15994 25764
rect 18049 25755 18107 25761
rect 18049 25721 18061 25755
rect 18095 25752 18107 25755
rect 18966 25752 18972 25764
rect 18095 25724 18972 25752
rect 18095 25721 18107 25724
rect 18049 25715 18107 25721
rect 18966 25712 18972 25724
rect 19024 25712 19030 25764
rect 1854 25644 1860 25696
rect 1912 25684 1918 25696
rect 2225 25687 2283 25693
rect 2225 25684 2237 25687
rect 1912 25656 2237 25684
rect 1912 25644 1918 25656
rect 2225 25653 2237 25656
rect 2271 25653 2283 25687
rect 2225 25647 2283 25653
rect 3513 25687 3571 25693
rect 3513 25653 3525 25687
rect 3559 25684 3571 25687
rect 3786 25684 3792 25696
rect 3559 25656 3792 25684
rect 3559 25653 3571 25656
rect 3513 25647 3571 25653
rect 3786 25644 3792 25656
rect 3844 25644 3850 25696
rect 3970 25644 3976 25696
rect 4028 25684 4034 25696
rect 4157 25687 4215 25693
rect 4157 25684 4169 25687
rect 4028 25656 4169 25684
rect 4028 25644 4034 25656
rect 4157 25653 4169 25656
rect 4203 25653 4215 25687
rect 4706 25684 4712 25696
rect 4667 25656 4712 25684
rect 4157 25647 4215 25653
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 8294 25684 8300 25696
rect 8255 25656 8300 25684
rect 8294 25644 8300 25656
rect 8352 25684 8358 25696
rect 10134 25684 10140 25696
rect 8352 25656 10140 25684
rect 8352 25644 8358 25656
rect 10134 25644 10140 25656
rect 10192 25644 10198 25696
rect 10226 25644 10232 25696
rect 10284 25684 10290 25696
rect 10873 25687 10931 25693
rect 10873 25684 10885 25687
rect 10284 25656 10885 25684
rect 10284 25644 10290 25656
rect 10873 25653 10885 25656
rect 10919 25653 10931 25687
rect 10873 25647 10931 25653
rect 11422 25644 11428 25696
rect 11480 25684 11486 25696
rect 12529 25687 12587 25693
rect 12529 25684 12541 25687
rect 11480 25656 12541 25684
rect 11480 25644 11486 25656
rect 12529 25653 12541 25656
rect 12575 25653 12587 25687
rect 12529 25647 12587 25653
rect 14090 25644 14096 25696
rect 14148 25684 14154 25696
rect 14185 25687 14243 25693
rect 14185 25684 14197 25687
rect 14148 25656 14197 25684
rect 14148 25644 14154 25656
rect 14185 25653 14197 25656
rect 14231 25653 14243 25687
rect 18782 25684 18788 25696
rect 18743 25656 18788 25684
rect 14185 25647 14243 25653
rect 18782 25644 18788 25656
rect 18840 25644 18846 25696
rect 19334 25684 19340 25696
rect 19295 25656 19340 25684
rect 19334 25644 19340 25656
rect 19392 25644 19398 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 5258 25480 5264 25492
rect 5219 25452 5264 25480
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 11882 25440 11888 25492
rect 11940 25480 11946 25492
rect 12805 25483 12863 25489
rect 12805 25480 12817 25483
rect 11940 25452 12817 25480
rect 11940 25440 11946 25452
rect 12805 25449 12817 25452
rect 12851 25449 12863 25483
rect 12805 25443 12863 25449
rect 12894 25440 12900 25492
rect 12952 25480 12958 25492
rect 17862 25480 17868 25492
rect 12952 25452 17868 25480
rect 12952 25440 12958 25452
rect 17862 25440 17868 25452
rect 17920 25440 17926 25492
rect 18782 25440 18788 25492
rect 18840 25480 18846 25492
rect 31110 25480 31116 25492
rect 18840 25452 31116 25480
rect 18840 25440 18846 25452
rect 31110 25440 31116 25452
rect 31168 25440 31174 25492
rect 32217 25483 32275 25489
rect 32217 25449 32229 25483
rect 32263 25480 32275 25483
rect 35894 25480 35900 25492
rect 32263 25452 35900 25480
rect 32263 25449 32275 25452
rect 32217 25443 32275 25449
rect 35894 25440 35900 25452
rect 35952 25440 35958 25492
rect 10778 25372 10784 25424
rect 10836 25412 10842 25424
rect 19705 25415 19763 25421
rect 10836 25384 18276 25412
rect 10836 25372 10842 25384
rect 12820 25356 12848 25384
rect 1857 25347 1915 25353
rect 1857 25313 1869 25347
rect 1903 25344 1915 25347
rect 7926 25344 7932 25356
rect 1903 25316 7932 25344
rect 1903 25313 1915 25316
rect 1857 25307 1915 25313
rect 7926 25304 7932 25316
rect 7984 25304 7990 25356
rect 11330 25344 11336 25356
rect 11291 25316 11336 25344
rect 11330 25304 11336 25316
rect 11388 25304 11394 25356
rect 12526 25304 12532 25356
rect 12584 25344 12590 25356
rect 12621 25347 12679 25353
rect 12621 25344 12633 25347
rect 12584 25316 12633 25344
rect 12584 25304 12590 25316
rect 12621 25313 12633 25316
rect 12667 25313 12679 25347
rect 12621 25307 12679 25313
rect 12802 25304 12808 25356
rect 12860 25304 12866 25356
rect 14918 25304 14924 25356
rect 14976 25344 14982 25356
rect 17126 25344 17132 25356
rect 14976 25316 17132 25344
rect 14976 25304 14982 25316
rect 17126 25304 17132 25316
rect 17184 25304 17190 25356
rect 17494 25344 17500 25356
rect 17455 25316 17500 25344
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 2869 25279 2927 25285
rect 2869 25276 2881 25279
rect 2746 25248 2881 25276
rect 1026 25168 1032 25220
rect 1084 25208 1090 25220
rect 2746 25208 2774 25248
rect 2869 25245 2881 25248
rect 2915 25245 2927 25279
rect 3970 25276 3976 25288
rect 3931 25248 3976 25276
rect 2869 25239 2927 25245
rect 3970 25236 3976 25248
rect 4028 25236 4034 25288
rect 4522 25236 4528 25288
rect 4580 25276 4586 25288
rect 4617 25279 4675 25285
rect 4617 25276 4629 25279
rect 4580 25248 4629 25276
rect 4580 25236 4586 25248
rect 4617 25245 4629 25248
rect 4663 25245 4675 25279
rect 4617 25239 4675 25245
rect 5350 25236 5356 25288
rect 5408 25276 5414 25288
rect 5445 25279 5503 25285
rect 5445 25276 5457 25279
rect 5408 25248 5457 25276
rect 5408 25236 5414 25248
rect 5445 25245 5457 25248
rect 5491 25245 5503 25279
rect 5445 25239 5503 25245
rect 8478 25236 8484 25288
rect 8536 25276 8542 25288
rect 9214 25276 9220 25288
rect 8536 25248 9220 25276
rect 8536 25236 8542 25248
rect 9214 25236 9220 25248
rect 9272 25276 9278 25288
rect 9585 25279 9643 25285
rect 9585 25276 9597 25279
rect 9272 25248 9597 25276
rect 9272 25236 9278 25248
rect 9585 25245 9597 25248
rect 9631 25245 9643 25279
rect 9585 25239 9643 25245
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25276 10471 25279
rect 12437 25279 12495 25285
rect 10459 25248 11192 25276
rect 10459 25245 10471 25248
rect 10413 25239 10471 25245
rect 1084 25180 2774 25208
rect 4065 25211 4123 25217
rect 1084 25168 1090 25180
rect 4065 25177 4077 25211
rect 4111 25208 4123 25211
rect 10778 25208 10784 25220
rect 4111 25180 10784 25208
rect 4111 25177 4123 25180
rect 4065 25171 4123 25177
rect 10778 25168 10784 25180
rect 10836 25168 10842 25220
rect 2961 25143 3019 25149
rect 2961 25109 2973 25143
rect 3007 25140 3019 25143
rect 3234 25140 3240 25152
rect 3007 25112 3240 25140
rect 3007 25109 3019 25112
rect 2961 25103 3019 25109
rect 3234 25100 3240 25112
rect 3292 25100 3298 25152
rect 4614 25100 4620 25152
rect 4672 25140 4678 25152
rect 4709 25143 4767 25149
rect 4709 25140 4721 25143
rect 4672 25112 4721 25140
rect 4672 25100 4678 25112
rect 4709 25109 4721 25112
rect 4755 25109 4767 25143
rect 4709 25103 4767 25109
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 6825 25143 6883 25149
rect 6825 25140 6837 25143
rect 6788 25112 6837 25140
rect 6788 25100 6794 25112
rect 6825 25109 6837 25112
rect 6871 25109 6883 25143
rect 9674 25140 9680 25152
rect 9635 25112 9680 25140
rect 6825 25103 6883 25109
rect 9674 25100 9680 25112
rect 9732 25100 9738 25152
rect 10134 25100 10140 25152
rect 10192 25140 10198 25152
rect 10505 25143 10563 25149
rect 10505 25140 10517 25143
rect 10192 25112 10517 25140
rect 10192 25100 10198 25112
rect 10505 25109 10517 25112
rect 10551 25109 10563 25143
rect 11164 25140 11192 25248
rect 12437 25245 12449 25279
rect 12483 25276 12495 25279
rect 13722 25276 13728 25288
rect 12483 25248 13728 25276
rect 12483 25245 12495 25248
rect 12437 25239 12495 25245
rect 13722 25236 13728 25248
rect 13780 25236 13786 25288
rect 18248 25285 18276 25384
rect 19705 25381 19717 25415
rect 19751 25412 19763 25415
rect 19978 25412 19984 25424
rect 19751 25384 19984 25412
rect 19751 25381 19763 25384
rect 19705 25375 19763 25381
rect 19978 25372 19984 25384
rect 20036 25372 20042 25424
rect 21545 25347 21603 25353
rect 21545 25313 21557 25347
rect 21591 25344 21603 25347
rect 22830 25344 22836 25356
rect 21591 25316 22836 25344
rect 21591 25313 21603 25316
rect 21545 25307 21603 25313
rect 22830 25304 22836 25316
rect 22888 25304 22894 25356
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25276 18291 25279
rect 18414 25276 18420 25288
rect 18279 25248 18420 25276
rect 18279 25245 18291 25248
rect 18233 25239 18291 25245
rect 18414 25236 18420 25248
rect 18472 25236 18478 25288
rect 19242 25236 19248 25288
rect 19300 25276 19306 25288
rect 19521 25279 19579 25285
rect 19521 25276 19533 25279
rect 19300 25248 19533 25276
rect 19300 25236 19306 25248
rect 19521 25245 19533 25248
rect 19567 25245 19579 25279
rect 19521 25239 19579 25245
rect 20717 25279 20775 25285
rect 20717 25245 20729 25279
rect 20763 25276 20775 25279
rect 21361 25279 21419 25285
rect 21361 25276 21373 25279
rect 20763 25248 21373 25276
rect 20763 25245 20775 25248
rect 20717 25239 20775 25245
rect 21361 25245 21373 25248
rect 21407 25245 21419 25279
rect 21361 25239 21419 25245
rect 24118 25236 24124 25288
rect 24176 25276 24182 25288
rect 27249 25279 27307 25285
rect 27249 25276 27261 25279
rect 24176 25248 27261 25276
rect 24176 25236 24182 25248
rect 27249 25245 27261 25248
rect 27295 25245 27307 25279
rect 27249 25239 27307 25245
rect 27341 25279 27399 25285
rect 27341 25245 27353 25279
rect 27387 25276 27399 25279
rect 32401 25279 32459 25285
rect 32401 25276 32413 25279
rect 27387 25248 32413 25276
rect 27387 25245 27399 25248
rect 27341 25239 27399 25245
rect 32401 25245 32413 25248
rect 32447 25245 32459 25279
rect 32401 25239 32459 25245
rect 11422 25168 11428 25220
rect 11480 25208 11486 25220
rect 11977 25211 12035 25217
rect 11480 25180 11525 25208
rect 11480 25168 11486 25180
rect 11977 25177 11989 25211
rect 12023 25208 12035 25211
rect 12066 25208 12072 25220
rect 12023 25180 12072 25208
rect 12023 25177 12035 25180
rect 11977 25171 12035 25177
rect 12066 25168 12072 25180
rect 12124 25168 12130 25220
rect 17221 25211 17279 25217
rect 17221 25177 17233 25211
rect 17267 25177 17279 25211
rect 17221 25171 17279 25177
rect 12894 25140 12900 25152
rect 11164 25112 12900 25140
rect 10505 25103 10563 25109
rect 12894 25100 12900 25112
rect 12952 25100 12958 25152
rect 16393 25143 16451 25149
rect 16393 25109 16405 25143
rect 16439 25140 16451 25143
rect 16942 25140 16948 25152
rect 16439 25112 16948 25140
rect 16439 25109 16451 25112
rect 16393 25103 16451 25109
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 17236 25140 17264 25171
rect 18325 25143 18383 25149
rect 18325 25140 18337 25143
rect 17236 25112 18337 25140
rect 18325 25109 18337 25112
rect 18371 25109 18383 25143
rect 18325 25103 18383 25109
rect 21910 25100 21916 25152
rect 21968 25140 21974 25152
rect 22005 25143 22063 25149
rect 22005 25140 22017 25143
rect 21968 25112 22017 25140
rect 21968 25100 21974 25112
rect 22005 25109 22017 25112
rect 22051 25109 22063 25143
rect 22005 25103 22063 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 6564 24908 6868 24936
rect 1946 24828 1952 24880
rect 2004 24868 2010 24880
rect 2498 24868 2504 24880
rect 2004 24840 2504 24868
rect 2004 24828 2010 24840
rect 2498 24828 2504 24840
rect 2556 24828 2562 24880
rect 5626 24868 5632 24880
rect 3620 24840 3924 24868
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24769 2283 24803
rect 2682 24800 2688 24812
rect 2643 24772 2688 24800
rect 2225 24763 2283 24769
rect 2240 24732 2268 24763
rect 2682 24760 2688 24772
rect 2740 24760 2746 24812
rect 3418 24760 3424 24812
rect 3476 24800 3482 24812
rect 3620 24800 3648 24840
rect 3476 24772 3648 24800
rect 3476 24760 3482 24772
rect 3694 24760 3700 24812
rect 3752 24800 3758 24812
rect 3789 24803 3847 24809
rect 3789 24800 3801 24803
rect 3752 24772 3801 24800
rect 3752 24760 3758 24772
rect 3789 24769 3801 24772
rect 3835 24769 3847 24803
rect 3896 24800 3924 24840
rect 5092 24840 5632 24868
rect 4522 24800 4528 24812
rect 3896 24772 4528 24800
rect 3789 24763 3847 24769
rect 4522 24760 4528 24772
rect 4580 24800 4586 24812
rect 5092 24809 5120 24840
rect 5626 24828 5632 24840
rect 5684 24828 5690 24880
rect 6564 24812 6592 24908
rect 6730 24868 6736 24880
rect 6691 24840 6736 24868
rect 6730 24828 6736 24840
rect 6788 24828 6794 24880
rect 6840 24877 6868 24908
rect 12066 24896 12072 24948
rect 12124 24936 12130 24948
rect 17494 24936 17500 24948
rect 12124 24908 17500 24936
rect 12124 24896 12130 24908
rect 17494 24896 17500 24908
rect 17552 24936 17558 24948
rect 23569 24939 23627 24945
rect 17552 24908 17632 24936
rect 17552 24896 17558 24908
rect 6825 24871 6883 24877
rect 6825 24837 6837 24871
rect 6871 24837 6883 24871
rect 8110 24868 8116 24880
rect 8071 24840 8116 24868
rect 6825 24831 6883 24837
rect 8110 24828 8116 24840
rect 8168 24828 8174 24880
rect 9306 24868 9312 24880
rect 9267 24840 9312 24868
rect 9306 24828 9312 24840
rect 9364 24828 9370 24880
rect 14090 24868 14096 24880
rect 11716 24840 11928 24868
rect 14051 24840 14096 24868
rect 4617 24803 4675 24809
rect 4617 24800 4629 24803
rect 4580 24772 4629 24800
rect 4580 24760 4586 24772
rect 4617 24769 4629 24772
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 5077 24803 5135 24809
rect 5077 24769 5089 24803
rect 5123 24769 5135 24803
rect 5077 24763 5135 24769
rect 5534 24760 5540 24812
rect 5592 24800 5598 24812
rect 5905 24803 5963 24809
rect 5905 24800 5917 24803
rect 5592 24772 5917 24800
rect 5592 24760 5598 24772
rect 5905 24769 5917 24772
rect 5951 24769 5963 24803
rect 5905 24763 5963 24769
rect 6546 24760 6552 24812
rect 6604 24760 6610 24812
rect 10962 24760 10968 24812
rect 11020 24800 11026 24812
rect 11716 24800 11744 24840
rect 11020 24772 11744 24800
rect 11793 24803 11851 24809
rect 11020 24760 11026 24772
rect 11793 24769 11805 24803
rect 11839 24769 11851 24803
rect 11793 24763 11851 24769
rect 6178 24732 6184 24744
rect 2240 24704 6184 24732
rect 6178 24692 6184 24704
rect 6236 24692 6242 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7944 24704 8033 24732
rect 7944 24676 7972 24704
rect 8021 24701 8033 24704
rect 8067 24701 8079 24735
rect 8021 24695 8079 24701
rect 8202 24692 8208 24744
rect 8260 24732 8266 24744
rect 8297 24735 8355 24741
rect 8297 24732 8309 24735
rect 8260 24704 8309 24732
rect 8260 24692 8266 24704
rect 8297 24701 8309 24704
rect 8343 24701 8355 24735
rect 9214 24732 9220 24744
rect 9175 24704 9220 24732
rect 8297 24695 8355 24701
rect 9214 24692 9220 24704
rect 9272 24692 9278 24744
rect 9398 24692 9404 24744
rect 9456 24732 9462 24744
rect 11808 24732 11836 24763
rect 9456 24704 11836 24732
rect 11900 24732 11928 24840
rect 14090 24828 14096 24840
rect 14148 24828 14154 24880
rect 17604 24877 17632 24908
rect 23569 24905 23581 24939
rect 23615 24936 23627 24939
rect 23615 24908 23888 24936
rect 23615 24905 23627 24908
rect 23569 24899 23627 24905
rect 17037 24871 17095 24877
rect 17037 24868 17049 24871
rect 16776 24840 17049 24868
rect 13265 24803 13323 24809
rect 13265 24769 13277 24803
rect 13311 24800 13323 24803
rect 13814 24800 13820 24812
rect 13311 24772 13820 24800
rect 13311 24769 13323 24772
rect 13265 24763 13323 24769
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 15102 24800 15108 24812
rect 14844 24772 15108 24800
rect 14001 24735 14059 24741
rect 11900 24704 13952 24732
rect 9456 24692 9462 24704
rect 5721 24667 5779 24673
rect 5721 24664 5733 24667
rect 3712 24636 5733 24664
rect 2038 24596 2044 24608
rect 1999 24568 2044 24596
rect 2038 24556 2044 24568
rect 2096 24556 2102 24608
rect 2774 24556 2780 24608
rect 2832 24596 2838 24608
rect 2832 24568 2877 24596
rect 2832 24556 2838 24568
rect 3050 24556 3056 24608
rect 3108 24596 3114 24608
rect 3712 24596 3740 24636
rect 5721 24633 5733 24636
rect 5767 24633 5779 24667
rect 5721 24627 5779 24633
rect 7285 24667 7343 24673
rect 7285 24633 7297 24667
rect 7331 24633 7343 24667
rect 7285 24627 7343 24633
rect 3878 24596 3884 24608
rect 3108 24568 3740 24596
rect 3839 24568 3884 24596
rect 3108 24556 3114 24568
rect 3878 24556 3884 24568
rect 3936 24556 3942 24608
rect 4433 24599 4491 24605
rect 4433 24565 4445 24599
rect 4479 24596 4491 24599
rect 4982 24596 4988 24608
rect 4479 24568 4988 24596
rect 4479 24565 4491 24568
rect 4433 24559 4491 24565
rect 4982 24556 4988 24568
rect 5040 24556 5046 24608
rect 5169 24599 5227 24605
rect 5169 24565 5181 24599
rect 5215 24596 5227 24599
rect 5258 24596 5264 24608
rect 5215 24568 5264 24596
rect 5215 24565 5227 24568
rect 5169 24559 5227 24565
rect 5258 24556 5264 24568
rect 5316 24556 5322 24608
rect 7300 24596 7328 24627
rect 7926 24624 7932 24676
rect 7984 24624 7990 24676
rect 7558 24596 7564 24608
rect 7300 24568 7564 24596
rect 7558 24556 7564 24568
rect 7616 24596 7622 24608
rect 8220 24596 8248 24692
rect 8938 24624 8944 24676
rect 8996 24664 9002 24676
rect 9769 24667 9827 24673
rect 9769 24664 9781 24667
rect 8996 24636 9781 24664
rect 8996 24624 9002 24636
rect 9769 24633 9781 24636
rect 9815 24633 9827 24667
rect 9769 24627 9827 24633
rect 11698 24624 11704 24676
rect 11756 24664 11762 24676
rect 13170 24664 13176 24676
rect 11756 24636 13176 24664
rect 11756 24624 11762 24636
rect 13170 24624 13176 24636
rect 13228 24624 13234 24676
rect 13924 24664 13952 24704
rect 14001 24701 14013 24735
rect 14047 24732 14059 24735
rect 14366 24732 14372 24744
rect 14047 24704 14372 24732
rect 14047 24701 14059 24704
rect 14001 24695 14059 24701
rect 14366 24692 14372 24704
rect 14424 24692 14430 24744
rect 14844 24732 14872 24772
rect 15102 24760 15108 24772
rect 15160 24760 15166 24812
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 16117 24763 16175 24769
rect 16209 24803 16267 24809
rect 16209 24769 16221 24803
rect 16255 24800 16267 24803
rect 16776 24800 16804 24840
rect 17037 24837 17049 24840
rect 17083 24837 17095 24871
rect 17037 24831 17095 24837
rect 17589 24871 17647 24877
rect 17589 24837 17601 24871
rect 17635 24837 17647 24871
rect 22186 24868 22192 24880
rect 22147 24840 22192 24868
rect 17589 24831 17647 24837
rect 22186 24828 22192 24840
rect 22244 24828 22250 24880
rect 16255 24772 16804 24800
rect 18049 24803 18107 24809
rect 16255 24769 16267 24772
rect 16209 24763 16267 24769
rect 18049 24769 18061 24803
rect 18095 24800 18107 24803
rect 18138 24800 18144 24812
rect 18095 24772 18144 24800
rect 18095 24769 18107 24772
rect 18049 24763 18107 24769
rect 14476 24704 14872 24732
rect 16132 24732 16160 24763
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 18233 24803 18291 24809
rect 18233 24769 18245 24803
rect 18279 24800 18291 24803
rect 19334 24800 19340 24812
rect 18279 24772 19340 24800
rect 18279 24769 18291 24772
rect 18233 24763 18291 24769
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 20162 24800 20168 24812
rect 20123 24772 20168 24800
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 22830 24760 22836 24812
rect 22888 24800 22894 24812
rect 23753 24803 23811 24809
rect 23753 24800 23765 24803
rect 22888 24772 23765 24800
rect 22888 24760 22894 24772
rect 23753 24769 23765 24772
rect 23799 24769 23811 24803
rect 23860 24800 23888 24908
rect 24397 24803 24455 24809
rect 24397 24800 24409 24803
rect 23860 24772 24409 24800
rect 23753 24763 23811 24769
rect 24397 24769 24409 24772
rect 24443 24769 24455 24803
rect 24397 24763 24455 24769
rect 28997 24803 29055 24809
rect 28997 24769 29009 24803
rect 29043 24800 29055 24803
rect 29043 24772 31754 24800
rect 29043 24769 29055 24772
rect 28997 24763 29055 24769
rect 16942 24732 16948 24744
rect 16132 24704 16252 24732
rect 16903 24704 16948 24732
rect 14476 24664 14504 24704
rect 16224 24676 16252 24704
rect 16942 24692 16948 24704
rect 17000 24692 17006 24744
rect 19426 24692 19432 24744
rect 19484 24732 19490 24744
rect 19981 24735 20039 24741
rect 19981 24732 19993 24735
rect 19484 24704 19993 24732
rect 19484 24692 19490 24704
rect 19981 24701 19993 24704
rect 20027 24701 20039 24735
rect 19981 24695 20039 24701
rect 20625 24735 20683 24741
rect 20625 24701 20637 24735
rect 20671 24732 20683 24735
rect 21910 24732 21916 24744
rect 20671 24704 21916 24732
rect 20671 24701 20683 24704
rect 20625 24695 20683 24701
rect 21910 24692 21916 24704
rect 21968 24732 21974 24744
rect 22097 24735 22155 24741
rect 22097 24732 22109 24735
rect 21968 24704 22109 24732
rect 21968 24692 21974 24704
rect 22097 24701 22109 24704
rect 22143 24701 22155 24735
rect 31726 24732 31754 24772
rect 34514 24760 34520 24812
rect 34572 24800 34578 24812
rect 38013 24803 38071 24809
rect 38013 24800 38025 24803
rect 34572 24772 38025 24800
rect 34572 24760 34578 24772
rect 38013 24769 38025 24772
rect 38059 24769 38071 24803
rect 38013 24763 38071 24769
rect 35986 24732 35992 24744
rect 31726 24704 35992 24732
rect 22097 24695 22155 24701
rect 35986 24692 35992 24704
rect 36044 24692 36050 24744
rect 13924 24636 14504 24664
rect 14553 24667 14611 24673
rect 14553 24633 14565 24667
rect 14599 24633 14611 24667
rect 14553 24627 14611 24633
rect 11882 24596 11888 24608
rect 7616 24568 8248 24596
rect 11843 24568 11888 24596
rect 7616 24556 7622 24568
rect 11882 24556 11888 24568
rect 11940 24556 11946 24608
rect 13354 24596 13360 24608
rect 13315 24568 13360 24596
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 14568 24596 14596 24627
rect 14642 24624 14648 24676
rect 14700 24664 14706 24676
rect 16206 24664 16212 24676
rect 14700 24636 16068 24664
rect 16119 24636 16212 24664
rect 14700 24624 14706 24636
rect 15194 24596 15200 24608
rect 13596 24568 14596 24596
rect 15155 24568 15200 24596
rect 13596 24556 13602 24568
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 16040 24596 16068 24636
rect 16206 24624 16212 24636
rect 16264 24664 16270 24676
rect 20162 24664 20168 24676
rect 16264 24636 20168 24664
rect 16264 24624 16270 24636
rect 20162 24624 20168 24636
rect 20220 24624 20226 24676
rect 20898 24624 20904 24676
rect 20956 24664 20962 24676
rect 22649 24667 22707 24673
rect 22649 24664 22661 24667
rect 20956 24636 22661 24664
rect 20956 24624 20962 24636
rect 22649 24633 22661 24636
rect 22695 24664 22707 24667
rect 26234 24664 26240 24676
rect 22695 24636 26240 24664
rect 22695 24633 22707 24636
rect 22649 24627 22707 24633
rect 26234 24624 26240 24636
rect 26292 24624 26298 24676
rect 17034 24596 17040 24608
rect 16040 24568 17040 24596
rect 17034 24556 17040 24568
rect 17092 24556 17098 24608
rect 18690 24596 18696 24608
rect 18651 24568 18696 24596
rect 18690 24556 18696 24568
rect 18748 24556 18754 24608
rect 22186 24556 22192 24608
rect 22244 24596 22250 24608
rect 24213 24599 24271 24605
rect 24213 24596 24225 24599
rect 22244 24568 24225 24596
rect 22244 24556 22250 24568
rect 24213 24565 24225 24568
rect 24259 24565 24271 24599
rect 29086 24596 29092 24608
rect 29047 24568 29092 24596
rect 24213 24559 24271 24565
rect 29086 24556 29092 24568
rect 29144 24556 29150 24608
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 934 24352 940 24404
rect 992 24392 998 24404
rect 3694 24392 3700 24404
rect 992 24364 3700 24392
rect 992 24352 998 24364
rect 3694 24352 3700 24364
rect 3752 24352 3758 24404
rect 6178 24392 6184 24404
rect 6139 24364 6184 24392
rect 6178 24352 6184 24364
rect 6236 24352 6242 24404
rect 7834 24352 7840 24404
rect 7892 24392 7898 24404
rect 10502 24392 10508 24404
rect 7892 24364 10508 24392
rect 7892 24352 7898 24364
rect 10502 24352 10508 24364
rect 10560 24352 10566 24404
rect 11882 24352 11888 24404
rect 11940 24392 11946 24404
rect 13078 24392 13084 24404
rect 11940 24364 13084 24392
rect 11940 24352 11946 24364
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 13170 24352 13176 24404
rect 13228 24392 13234 24404
rect 16206 24392 16212 24404
rect 13228 24364 16212 24392
rect 13228 24352 13234 24364
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 17770 24352 17776 24404
rect 17828 24352 17834 24404
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 23569 24395 23627 24401
rect 23569 24392 23581 24395
rect 20128 24364 23581 24392
rect 20128 24352 20134 24364
rect 23569 24361 23581 24364
rect 23615 24361 23627 24395
rect 23569 24355 23627 24361
rect 3878 24284 3884 24336
rect 3936 24324 3942 24336
rect 12710 24324 12716 24336
rect 3936 24296 12716 24324
rect 3936 24284 3942 24296
rect 12710 24284 12716 24296
rect 12768 24284 12774 24336
rect 13262 24324 13268 24336
rect 13004 24296 13268 24324
rect 4338 24216 4344 24268
rect 4396 24256 4402 24268
rect 8021 24259 8079 24265
rect 4396 24228 7972 24256
rect 4396 24216 4402 24228
rect 1486 24148 1492 24200
rect 1544 24188 1550 24200
rect 1857 24191 1915 24197
rect 1857 24188 1869 24191
rect 1544 24160 1869 24188
rect 1544 24148 1550 24160
rect 1857 24157 1869 24160
rect 1903 24157 1915 24191
rect 2498 24188 2504 24200
rect 2459 24160 2504 24188
rect 1857 24151 1915 24157
rect 2498 24148 2504 24160
rect 2556 24148 2562 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4706 24188 4712 24200
rect 4203 24160 4712 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 4982 24188 4988 24200
rect 4943 24160 4988 24188
rect 4982 24148 4988 24160
rect 5040 24148 5046 24200
rect 5445 24191 5503 24197
rect 5445 24157 5457 24191
rect 5491 24188 5503 24191
rect 5626 24188 5632 24200
rect 5491 24160 5632 24188
rect 5491 24157 5503 24160
rect 5445 24151 5503 24157
rect 5626 24148 5632 24160
rect 5684 24148 5690 24200
rect 6086 24188 6092 24200
rect 6047 24160 6092 24188
rect 6086 24148 6092 24160
rect 6144 24148 6150 24200
rect 7009 24191 7067 24197
rect 7009 24157 7021 24191
rect 7055 24188 7067 24191
rect 7944 24188 7972 24228
rect 8021 24225 8033 24259
rect 8067 24256 8079 24259
rect 9214 24256 9220 24268
rect 8067 24228 9220 24256
rect 8067 24225 8079 24228
rect 8021 24219 8079 24225
rect 9214 24216 9220 24228
rect 9272 24216 9278 24268
rect 12526 24216 12532 24268
rect 12584 24256 12590 24268
rect 13004 24256 13032 24296
rect 13262 24284 13268 24296
rect 13320 24284 13326 24336
rect 17788 24324 17816 24352
rect 13740 24296 17816 24324
rect 13170 24256 13176 24268
rect 12584 24228 13032 24256
rect 13083 24228 13176 24256
rect 12584 24216 12590 24228
rect 13170 24216 13176 24228
rect 13228 24256 13234 24268
rect 13538 24256 13544 24268
rect 13228 24228 13544 24256
rect 13228 24216 13234 24228
rect 13538 24216 13544 24228
rect 13596 24216 13602 24268
rect 8294 24188 8300 24200
rect 7055 24160 7880 24188
rect 7944 24160 8300 24188
rect 7055 24157 7067 24160
rect 7009 24151 7067 24157
rect 2593 24123 2651 24129
rect 2593 24089 2605 24123
rect 2639 24120 2651 24123
rect 3602 24120 3608 24132
rect 2639 24092 3608 24120
rect 2639 24089 2651 24092
rect 2593 24083 2651 24089
rect 3602 24080 3608 24092
rect 3660 24080 3666 24132
rect 1949 24055 2007 24061
rect 1949 24021 1961 24055
rect 1995 24052 2007 24055
rect 2498 24052 2504 24064
rect 1995 24024 2504 24052
rect 1995 24021 2007 24024
rect 1949 24015 2007 24021
rect 2498 24012 2504 24024
rect 2556 24012 2562 24064
rect 3142 24052 3148 24064
rect 3103 24024 3148 24052
rect 3142 24012 3148 24024
rect 3200 24012 3206 24064
rect 3326 24012 3332 24064
rect 3384 24052 3390 24064
rect 4249 24055 4307 24061
rect 4249 24052 4261 24055
rect 3384 24024 4261 24052
rect 3384 24012 3390 24024
rect 4249 24021 4261 24024
rect 4295 24021 4307 24055
rect 4249 24015 4307 24021
rect 4706 24012 4712 24064
rect 4764 24052 4770 24064
rect 4801 24055 4859 24061
rect 4801 24052 4813 24055
rect 4764 24024 4813 24052
rect 4764 24012 4770 24024
rect 4801 24021 4813 24024
rect 4847 24021 4859 24055
rect 4801 24015 4859 24021
rect 4982 24012 4988 24064
rect 5040 24052 5046 24064
rect 5537 24055 5595 24061
rect 5537 24052 5549 24055
rect 5040 24024 5549 24052
rect 5040 24012 5046 24024
rect 5537 24021 5549 24024
rect 5583 24021 5595 24055
rect 7098 24052 7104 24064
rect 7059 24024 7104 24052
rect 5537 24015 5595 24021
rect 7098 24012 7104 24024
rect 7156 24012 7162 24064
rect 7852 24052 7880 24160
rect 8294 24148 8300 24160
rect 8352 24148 8358 24200
rect 10962 24148 10968 24200
rect 11020 24188 11026 24200
rect 11149 24191 11207 24197
rect 11149 24188 11161 24191
rect 11020 24160 11161 24188
rect 11020 24148 11026 24160
rect 11149 24157 11161 24160
rect 11195 24157 11207 24191
rect 13740 24188 13768 24296
rect 18046 24284 18052 24336
rect 18104 24324 18110 24336
rect 20898 24324 20904 24336
rect 18104 24296 20484 24324
rect 20859 24296 20904 24324
rect 18104 24284 18110 24296
rect 13814 24216 13820 24268
rect 13872 24256 13878 24268
rect 17770 24256 17776 24268
rect 13872 24228 17776 24256
rect 13872 24216 13878 24228
rect 14292 24197 14320 24228
rect 17770 24216 17776 24228
rect 17828 24216 17834 24268
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 17920 24228 18184 24256
rect 17920 24216 17926 24228
rect 11149 24151 11207 24157
rect 13188 24160 13768 24188
rect 14277 24191 14335 24197
rect 9122 24080 9128 24132
rect 9180 24120 9186 24132
rect 10045 24123 10103 24129
rect 10045 24120 10057 24123
rect 9180 24092 10057 24120
rect 9180 24080 9186 24092
rect 10045 24089 10057 24092
rect 10091 24089 10103 24123
rect 10045 24083 10103 24089
rect 10137 24123 10195 24129
rect 10137 24089 10149 24123
rect 10183 24120 10195 24123
rect 10226 24120 10232 24132
rect 10183 24092 10232 24120
rect 10183 24089 10195 24092
rect 10137 24083 10195 24089
rect 10226 24080 10232 24092
rect 10284 24080 10290 24132
rect 10686 24120 10692 24132
rect 10647 24092 10692 24120
rect 10686 24080 10692 24092
rect 10744 24080 10750 24132
rect 12618 24080 12624 24132
rect 12676 24120 12682 24132
rect 12676 24092 12721 24120
rect 12676 24080 12682 24092
rect 12986 24080 12992 24132
rect 13044 24120 13050 24132
rect 13188 24120 13216 24160
rect 14277 24157 14289 24191
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 14921 24191 14979 24197
rect 14921 24157 14933 24191
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 14936 24120 14964 24151
rect 15102 24148 15108 24200
rect 15160 24188 15166 24200
rect 18156 24197 18184 24228
rect 18690 24216 18696 24268
rect 18748 24256 18754 24268
rect 20349 24259 20407 24265
rect 20349 24256 20361 24259
rect 18748 24228 20361 24256
rect 18748 24216 18754 24228
rect 20349 24225 20361 24228
rect 20395 24225 20407 24259
rect 20456 24256 20484 24296
rect 20898 24284 20904 24296
rect 20956 24284 20962 24336
rect 20456 24228 22094 24256
rect 20349 24219 20407 24225
rect 16853 24191 16911 24197
rect 16853 24190 16865 24191
rect 16776 24188 16865 24190
rect 15160 24162 16865 24188
rect 15160 24160 16804 24162
rect 15160 24148 15166 24160
rect 16853 24157 16865 24162
rect 16899 24157 16911 24191
rect 16853 24151 16911 24157
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 18322 24148 18328 24200
rect 18380 24188 18386 24200
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 18380 24160 19441 24188
rect 18380 24148 18386 24160
rect 19429 24157 19441 24160
rect 19475 24188 19487 24191
rect 19518 24188 19524 24200
rect 19475 24160 19524 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 22066 24188 22094 24228
rect 22830 24188 22836 24200
rect 22066 24160 22836 24188
rect 22830 24148 22836 24160
rect 22888 24148 22894 24200
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24188 23811 24191
rect 24302 24188 24308 24200
rect 23799 24160 24308 24188
rect 23799 24157 23811 24160
rect 23753 24151 23811 24157
rect 24302 24148 24308 24160
rect 24360 24148 24366 24200
rect 36078 24148 36084 24200
rect 36136 24188 36142 24200
rect 38013 24191 38071 24197
rect 38013 24188 38025 24191
rect 36136 24160 38025 24188
rect 36136 24148 36142 24160
rect 38013 24157 38025 24160
rect 38059 24157 38071 24191
rect 38013 24151 38071 24157
rect 13044 24092 13216 24120
rect 13280 24092 14964 24120
rect 18233 24123 18291 24129
rect 13044 24080 13050 24092
rect 9766 24052 9772 24064
rect 7852 24024 9772 24052
rect 9766 24012 9772 24024
rect 9824 24012 9830 24064
rect 11238 24052 11244 24064
rect 11199 24024 11244 24052
rect 11238 24012 11244 24024
rect 11296 24012 11302 24064
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 13280 24052 13308 24092
rect 18233 24089 18245 24123
rect 18279 24120 18291 24123
rect 19334 24120 19340 24132
rect 18279 24092 19340 24120
rect 18279 24089 18291 24092
rect 18233 24083 18291 24089
rect 19334 24080 19340 24092
rect 19392 24080 19398 24132
rect 20441 24123 20499 24129
rect 20441 24089 20453 24123
rect 20487 24089 20499 24123
rect 20441 24083 20499 24089
rect 14366 24052 14372 24064
rect 12492 24024 13308 24052
rect 14327 24024 14372 24052
rect 12492 24012 12498 24024
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 15010 24052 15016 24064
rect 14971 24024 15016 24052
rect 15010 24012 15016 24024
rect 15068 24012 15074 24064
rect 16945 24055 17003 24061
rect 16945 24021 16957 24055
rect 16991 24052 17003 24055
rect 17586 24052 17592 24064
rect 16991 24024 17592 24052
rect 16991 24021 17003 24024
rect 16945 24015 17003 24021
rect 17586 24012 17592 24024
rect 17644 24012 17650 24064
rect 19242 24012 19248 24064
rect 19300 24052 19306 24064
rect 19521 24055 19579 24061
rect 19521 24052 19533 24055
rect 19300 24024 19533 24052
rect 19300 24012 19306 24024
rect 19521 24021 19533 24024
rect 19567 24021 19579 24055
rect 20456 24052 20484 24083
rect 22925 24055 22983 24061
rect 22925 24052 22937 24055
rect 20456 24024 22937 24052
rect 19521 24015 19579 24021
rect 22925 24021 22937 24024
rect 22971 24021 22983 24055
rect 38194 24052 38200 24064
rect 38155 24024 38200 24052
rect 22925 24015 22983 24021
rect 38194 24012 38200 24024
rect 38252 24012 38258 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 3602 23808 3608 23860
rect 3660 23848 3666 23860
rect 3660 23820 5304 23848
rect 3660 23808 3666 23820
rect 3329 23783 3387 23789
rect 3329 23749 3341 23783
rect 3375 23780 3387 23783
rect 4614 23780 4620 23792
rect 3375 23752 4620 23780
rect 3375 23749 3387 23752
rect 3329 23743 3387 23749
rect 4614 23740 4620 23752
rect 4672 23740 4678 23792
rect 5166 23780 5172 23792
rect 4908 23752 5172 23780
rect 1394 23672 1400 23724
rect 1452 23712 1458 23724
rect 1857 23715 1915 23721
rect 1857 23712 1869 23715
rect 1452 23684 1869 23712
rect 1452 23672 1458 23684
rect 1857 23681 1869 23684
rect 1903 23681 1915 23715
rect 1857 23675 1915 23681
rect 4341 23715 4399 23721
rect 4341 23681 4353 23715
rect 4387 23712 4399 23715
rect 4908 23712 4936 23752
rect 5166 23740 5172 23752
rect 5224 23740 5230 23792
rect 4387 23684 4936 23712
rect 4985 23715 5043 23721
rect 4387 23681 4399 23684
rect 4341 23675 4399 23681
rect 4985 23681 4997 23715
rect 5031 23681 5043 23715
rect 4985 23675 5043 23681
rect 2130 23644 2136 23656
rect 2091 23616 2136 23644
rect 2130 23604 2136 23616
rect 2188 23604 2194 23656
rect 3237 23647 3295 23653
rect 3237 23613 3249 23647
rect 3283 23613 3295 23647
rect 3237 23607 3295 23613
rect 1302 23536 1308 23588
rect 1360 23576 1366 23588
rect 3050 23576 3056 23588
rect 1360 23548 3056 23576
rect 1360 23536 1366 23548
rect 3050 23536 3056 23548
rect 3108 23536 3114 23588
rect 2038 23468 2044 23520
rect 2096 23508 2102 23520
rect 2682 23508 2688 23520
rect 2096 23480 2688 23508
rect 2096 23468 2102 23480
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 3252 23508 3280 23607
rect 3602 23604 3608 23656
rect 3660 23644 3666 23656
rect 5000 23644 5028 23675
rect 5074 23672 5080 23724
rect 5132 23712 5138 23724
rect 5276 23712 5304 23820
rect 5442 23808 5448 23860
rect 5500 23848 5506 23860
rect 7193 23851 7251 23857
rect 7193 23848 7205 23851
rect 5500 23820 7205 23848
rect 5500 23808 5506 23820
rect 7193 23817 7205 23820
rect 7239 23817 7251 23851
rect 9674 23848 9680 23860
rect 7193 23811 7251 23817
rect 8680 23820 9680 23848
rect 8570 23780 8576 23792
rect 8531 23752 8576 23780
rect 8570 23740 8576 23752
rect 8628 23740 8634 23792
rect 8680 23789 8708 23820
rect 9674 23808 9680 23820
rect 9732 23808 9738 23860
rect 10965 23851 11023 23857
rect 10965 23817 10977 23851
rect 11011 23817 11023 23851
rect 12434 23848 12440 23860
rect 10965 23811 11023 23817
rect 11808 23820 12440 23848
rect 8665 23783 8723 23789
rect 8665 23749 8677 23783
rect 8711 23749 8723 23783
rect 8665 23743 8723 23749
rect 5626 23712 5632 23724
rect 5132 23684 5304 23712
rect 5539 23684 5632 23712
rect 5132 23672 5138 23684
rect 5626 23672 5632 23684
rect 5684 23712 5690 23724
rect 6454 23712 6460 23724
rect 5684 23684 6460 23712
rect 5684 23672 5690 23684
rect 6454 23672 6460 23684
rect 6512 23712 6518 23724
rect 6549 23715 6607 23721
rect 6549 23712 6561 23715
rect 6512 23684 6561 23712
rect 6512 23672 6518 23684
rect 6549 23681 6561 23684
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 7006 23672 7012 23724
rect 7064 23712 7070 23724
rect 7377 23715 7435 23721
rect 7377 23712 7389 23715
rect 7064 23684 7389 23712
rect 7064 23672 7070 23684
rect 7377 23681 7389 23684
rect 7423 23681 7435 23715
rect 7834 23712 7840 23724
rect 7795 23684 7840 23712
rect 7377 23675 7435 23681
rect 7834 23672 7840 23684
rect 7892 23672 7898 23724
rect 9677 23715 9735 23721
rect 9677 23681 9689 23715
rect 9723 23712 9735 23715
rect 9766 23712 9772 23724
rect 9723 23684 9772 23712
rect 9723 23681 9735 23684
rect 9677 23675 9735 23681
rect 9766 23672 9772 23684
rect 9824 23712 9830 23724
rect 10318 23712 10324 23724
rect 9824 23684 10324 23712
rect 9824 23672 9830 23684
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23712 10563 23715
rect 10980 23712 11008 23811
rect 10551 23684 11008 23712
rect 10551 23681 10563 23684
rect 10505 23675 10563 23681
rect 11054 23672 11060 23724
rect 11112 23712 11118 23724
rect 11808 23721 11836 23820
rect 12434 23808 12440 23820
rect 12492 23808 12498 23860
rect 15010 23848 15016 23860
rect 12636 23820 15016 23848
rect 12636 23789 12664 23820
rect 15010 23808 15016 23820
rect 15068 23808 15074 23860
rect 15102 23808 15108 23860
rect 15160 23848 15166 23860
rect 18046 23848 18052 23860
rect 15160 23820 18052 23848
rect 15160 23808 15166 23820
rect 18046 23808 18052 23820
rect 18104 23808 18110 23860
rect 18690 23808 18696 23860
rect 18748 23848 18754 23860
rect 19705 23851 19763 23857
rect 19705 23848 19717 23851
rect 18748 23820 19717 23848
rect 18748 23808 18754 23820
rect 19705 23817 19717 23820
rect 19751 23817 19763 23851
rect 19705 23811 19763 23817
rect 19794 23808 19800 23860
rect 19852 23848 19858 23860
rect 29086 23848 29092 23860
rect 19852 23820 29092 23848
rect 19852 23808 19858 23820
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 12621 23783 12679 23789
rect 12621 23749 12633 23783
rect 12667 23749 12679 23783
rect 13722 23780 13728 23792
rect 13683 23752 13728 23780
rect 12621 23743 12679 23749
rect 13722 23740 13728 23752
rect 13780 23740 13786 23792
rect 13817 23783 13875 23789
rect 13817 23749 13829 23783
rect 13863 23780 13875 23783
rect 16025 23783 16083 23789
rect 16025 23780 16037 23783
rect 13863 23752 16037 23780
rect 13863 23749 13875 23752
rect 13817 23743 13875 23749
rect 16025 23749 16037 23752
rect 16071 23749 16083 23783
rect 17586 23780 17592 23792
rect 17547 23752 17592 23780
rect 16025 23743 16083 23749
rect 17586 23740 17592 23752
rect 17644 23740 17650 23792
rect 17770 23740 17776 23792
rect 17828 23780 17834 23792
rect 37734 23780 37740 23792
rect 17828 23752 37740 23780
rect 17828 23740 17834 23752
rect 37734 23740 37740 23752
rect 37792 23740 37798 23792
rect 11149 23715 11207 23721
rect 11149 23712 11161 23715
rect 11112 23684 11161 23712
rect 11112 23672 11118 23684
rect 11149 23681 11161 23684
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 11793 23715 11851 23721
rect 11793 23681 11805 23715
rect 11839 23681 11851 23715
rect 14826 23712 14832 23724
rect 14787 23684 14832 23712
rect 11793 23675 11851 23681
rect 5810 23644 5816 23656
rect 3660 23616 5028 23644
rect 5092 23616 5816 23644
rect 3660 23604 3666 23616
rect 3789 23579 3847 23585
rect 3789 23545 3801 23579
rect 3835 23576 3847 23579
rect 3970 23576 3976 23588
rect 3835 23548 3976 23576
rect 3835 23545 3847 23548
rect 3789 23539 3847 23545
rect 3970 23536 3976 23548
rect 4028 23576 4034 23588
rect 5092 23576 5120 23616
rect 5810 23604 5816 23616
rect 5868 23604 5874 23656
rect 6178 23604 6184 23656
rect 6236 23644 6242 23656
rect 7929 23647 7987 23653
rect 7929 23644 7941 23647
rect 6236 23616 7941 23644
rect 6236 23604 6242 23616
rect 7929 23613 7941 23616
rect 7975 23613 7987 23647
rect 11808 23644 11836 23675
rect 14826 23672 14832 23684
rect 14884 23672 14890 23724
rect 15930 23712 15936 23724
rect 15891 23684 15936 23712
rect 15930 23672 15936 23684
rect 15988 23672 15994 23724
rect 19242 23712 19248 23724
rect 19203 23684 19248 23712
rect 19242 23672 19248 23684
rect 19300 23672 19306 23724
rect 20162 23672 20168 23724
rect 20220 23712 20226 23724
rect 22557 23715 22615 23721
rect 22557 23712 22569 23715
rect 20220 23684 22569 23712
rect 20220 23672 20226 23684
rect 22557 23681 22569 23684
rect 22603 23681 22615 23715
rect 23474 23712 23480 23724
rect 23435 23684 23480 23712
rect 22557 23675 22615 23681
rect 7929 23607 7987 23613
rect 8036 23616 11836 23644
rect 12529 23647 12587 23653
rect 4028 23548 5120 23576
rect 4028 23536 4034 23548
rect 5994 23536 6000 23588
rect 6052 23576 6058 23588
rect 6641 23579 6699 23585
rect 6641 23576 6653 23579
rect 6052 23548 6653 23576
rect 6052 23536 6058 23548
rect 6641 23545 6653 23548
rect 6687 23545 6699 23579
rect 6641 23539 6699 23545
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 8036 23576 8064 23616
rect 12529 23613 12541 23647
rect 12575 23644 12587 23647
rect 12986 23644 12992 23656
rect 12575 23616 12992 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 12986 23604 12992 23616
rect 13044 23604 13050 23656
rect 13173 23647 13231 23653
rect 13173 23613 13185 23647
rect 13219 23613 13231 23647
rect 13173 23607 13231 23613
rect 7892 23548 8064 23576
rect 7892 23536 7898 23548
rect 8662 23536 8668 23588
rect 8720 23576 8726 23588
rect 9125 23579 9183 23585
rect 9125 23576 9137 23579
rect 8720 23548 9137 23576
rect 8720 23536 8726 23548
rect 9125 23545 9137 23548
rect 9171 23576 9183 23579
rect 13188 23576 13216 23607
rect 13722 23604 13728 23656
rect 13780 23644 13786 23656
rect 14921 23647 14979 23653
rect 14921 23644 14933 23647
rect 13780 23616 14933 23644
rect 13780 23604 13786 23616
rect 14921 23613 14933 23616
rect 14967 23613 14979 23647
rect 14921 23607 14979 23613
rect 17497 23647 17555 23653
rect 17497 23613 17509 23647
rect 17543 23613 17555 23647
rect 17954 23644 17960 23656
rect 17915 23616 17960 23644
rect 17497 23607 17555 23613
rect 13906 23576 13912 23588
rect 9171 23548 13912 23576
rect 9171 23545 9183 23548
rect 9125 23539 9183 23545
rect 13906 23536 13912 23548
rect 13964 23536 13970 23588
rect 14277 23579 14335 23585
rect 14277 23545 14289 23579
rect 14323 23576 14335 23579
rect 15654 23576 15660 23588
rect 14323 23548 15660 23576
rect 14323 23545 14335 23548
rect 14277 23539 14335 23545
rect 15654 23536 15660 23548
rect 15712 23536 15718 23588
rect 17512 23576 17540 23607
rect 17954 23604 17960 23616
rect 18012 23644 18018 23656
rect 18782 23644 18788 23656
rect 18012 23616 18788 23644
rect 18012 23604 18018 23616
rect 18782 23604 18788 23616
rect 18840 23604 18846 23656
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23644 19119 23647
rect 19518 23644 19524 23656
rect 19107 23616 19524 23644
rect 19107 23613 19119 23616
rect 19061 23607 19119 23613
rect 19518 23604 19524 23616
rect 19576 23644 19582 23656
rect 20346 23644 20352 23656
rect 19576 23616 20352 23644
rect 19576 23604 19582 23616
rect 20346 23604 20352 23616
rect 20404 23604 20410 23656
rect 22572 23644 22600 23675
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 31205 23715 31263 23721
rect 31205 23681 31217 23715
rect 31251 23712 31263 23715
rect 34606 23712 34612 23724
rect 31251 23684 34612 23712
rect 31251 23681 31263 23684
rect 31205 23675 31263 23681
rect 34606 23672 34612 23684
rect 34664 23672 34670 23724
rect 24578 23644 24584 23656
rect 22572 23616 24584 23644
rect 24578 23604 24584 23616
rect 24636 23604 24642 23656
rect 18230 23576 18236 23588
rect 17512 23548 18236 23576
rect 18230 23536 18236 23548
rect 18288 23536 18294 23588
rect 4338 23508 4344 23520
rect 3252 23480 4344 23508
rect 4338 23468 4344 23480
rect 4396 23468 4402 23520
rect 4433 23511 4491 23517
rect 4433 23477 4445 23511
rect 4479 23508 4491 23511
rect 4614 23508 4620 23520
rect 4479 23480 4620 23508
rect 4479 23477 4491 23480
rect 4433 23471 4491 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 5077 23511 5135 23517
rect 5077 23477 5089 23511
rect 5123 23508 5135 23511
rect 5166 23508 5172 23520
rect 5123 23480 5172 23508
rect 5123 23477 5135 23480
rect 5077 23471 5135 23477
rect 5166 23468 5172 23480
rect 5224 23468 5230 23520
rect 5626 23468 5632 23520
rect 5684 23508 5690 23520
rect 5721 23511 5779 23517
rect 5721 23508 5733 23511
rect 5684 23480 5733 23508
rect 5684 23468 5690 23480
rect 5721 23477 5733 23480
rect 5767 23477 5779 23511
rect 9766 23508 9772 23520
rect 9727 23480 9772 23508
rect 5721 23471 5779 23477
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 10321 23511 10379 23517
rect 10321 23477 10333 23511
rect 10367 23508 10379 23511
rect 10870 23508 10876 23520
rect 10367 23480 10876 23508
rect 10367 23477 10379 23480
rect 10321 23471 10379 23477
rect 10870 23468 10876 23480
rect 10928 23468 10934 23520
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12618 23508 12624 23520
rect 11931 23480 12624 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12618 23468 12624 23480
rect 12676 23468 12682 23520
rect 13078 23468 13084 23520
rect 13136 23508 13142 23520
rect 15470 23508 15476 23520
rect 13136 23480 15476 23508
rect 13136 23468 13142 23480
rect 15470 23468 15476 23480
rect 15528 23468 15534 23520
rect 17034 23468 17040 23520
rect 17092 23508 17098 23520
rect 19794 23508 19800 23520
rect 17092 23480 19800 23508
rect 17092 23468 17098 23480
rect 19794 23468 19800 23480
rect 19852 23468 19858 23520
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 22649 23511 22707 23517
rect 22649 23508 22661 23511
rect 20036 23480 22661 23508
rect 20036 23468 20042 23480
rect 22649 23477 22661 23480
rect 22695 23477 22707 23511
rect 23290 23508 23296 23520
rect 23251 23480 23296 23508
rect 22649 23471 22707 23477
rect 23290 23468 23296 23480
rect 23348 23468 23354 23520
rect 28994 23468 29000 23520
rect 29052 23508 29058 23520
rect 31297 23511 31355 23517
rect 31297 23508 31309 23511
rect 29052 23480 31309 23508
rect 29052 23468 29058 23480
rect 31297 23477 31309 23480
rect 31343 23477 31355 23511
rect 31297 23471 31355 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 3329 23307 3387 23313
rect 3329 23273 3341 23307
rect 3375 23304 3387 23307
rect 6546 23304 6552 23316
rect 3375 23276 6552 23304
rect 3375 23273 3387 23276
rect 3329 23267 3387 23273
rect 6546 23264 6552 23276
rect 6604 23264 6610 23316
rect 7926 23264 7932 23316
rect 7984 23304 7990 23316
rect 7984 23276 11468 23304
rect 7984 23264 7990 23276
rect 3510 23196 3516 23248
rect 3568 23236 3574 23248
rect 4798 23236 4804 23248
rect 3568 23208 4804 23236
rect 3568 23196 3574 23208
rect 4798 23196 4804 23208
rect 4856 23196 4862 23248
rect 8846 23236 8852 23248
rect 6564 23208 8852 23236
rect 2958 23168 2964 23180
rect 1596 23140 2964 23168
rect 1596 22964 1624 23140
rect 2958 23128 2964 23140
rect 3016 23128 3022 23180
rect 4157 23171 4215 23177
rect 4157 23137 4169 23171
rect 4203 23168 4215 23171
rect 6564 23168 6592 23208
rect 8846 23196 8852 23208
rect 8904 23196 8910 23248
rect 10520 23245 10548 23276
rect 10505 23239 10563 23245
rect 10505 23205 10517 23239
rect 10551 23205 10563 23239
rect 10505 23199 10563 23205
rect 4203 23140 6592 23168
rect 6656 23140 7972 23168
rect 4203 23137 4215 23140
rect 4157 23131 4215 23137
rect 3050 23060 3056 23112
rect 3108 23100 3114 23112
rect 3237 23103 3295 23109
rect 3237 23100 3249 23103
rect 3108 23072 3249 23100
rect 3108 23060 3114 23072
rect 3237 23069 3249 23072
rect 3283 23069 3295 23103
rect 4062 23100 4068 23112
rect 4023 23072 4068 23100
rect 3237 23063 3295 23069
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 4801 23103 4859 23109
rect 4801 23069 4813 23103
rect 4847 23100 4859 23103
rect 5718 23100 5724 23112
rect 4847 23072 5724 23100
rect 4847 23069 4859 23072
rect 4801 23063 4859 23069
rect 5718 23060 5724 23072
rect 5776 23060 5782 23112
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23100 5871 23103
rect 6362 23100 6368 23112
rect 5859 23072 6368 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 6362 23060 6368 23072
rect 6420 23060 6426 23112
rect 6457 23103 6515 23109
rect 6457 23069 6469 23103
rect 6503 23100 6515 23103
rect 6656 23100 6684 23140
rect 6503 23072 6684 23100
rect 6503 23069 6515 23072
rect 6457 23063 6515 23069
rect 1762 23032 1768 23044
rect 1723 23004 1768 23032
rect 1762 22992 1768 23004
rect 1820 22992 1826 23044
rect 1857 23035 1915 23041
rect 1857 23001 1869 23035
rect 1903 23001 1915 23035
rect 1857 22995 1915 23001
rect 2409 23035 2467 23041
rect 2409 23001 2421 23035
rect 2455 23032 2467 23035
rect 3786 23032 3792 23044
rect 2455 23004 3792 23032
rect 2455 23001 2467 23004
rect 2409 22995 2467 23001
rect 1872 22964 1900 22995
rect 3786 22992 3792 23004
rect 3844 22992 3850 23044
rect 6549 23035 6607 23041
rect 6549 23032 6561 23035
rect 5828 23004 6561 23032
rect 5828 22976 5856 23004
rect 6549 23001 6561 23004
rect 6595 23001 6607 23035
rect 6656 23032 6684 23072
rect 6822 23060 6828 23112
rect 6880 23100 6886 23112
rect 7944 23109 7972 23140
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 11146 23168 11152 23180
rect 9548 23140 10732 23168
rect 11107 23140 11152 23168
rect 9548 23128 9554 23140
rect 7101 23103 7159 23109
rect 7101 23100 7113 23103
rect 6880 23072 7113 23100
rect 6880 23060 6886 23072
rect 7101 23069 7113 23072
rect 7147 23069 7159 23103
rect 7101 23063 7159 23069
rect 7929 23103 7987 23109
rect 7929 23069 7941 23103
rect 7975 23069 7987 23103
rect 7929 23063 7987 23069
rect 8570 23060 8576 23112
rect 8628 23100 8634 23112
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 8628 23072 9229 23100
rect 8628 23060 8634 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 6914 23032 6920 23044
rect 6656 23004 6920 23032
rect 6549 22995 6607 23001
rect 6914 22992 6920 23004
rect 6972 22992 6978 23044
rect 9674 23032 9680 23044
rect 7116 23004 9680 23032
rect 1596 22936 1900 22964
rect 2590 22924 2596 22976
rect 2648 22964 2654 22976
rect 3510 22964 3516 22976
rect 2648 22936 3516 22964
rect 2648 22924 2654 22936
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 4893 22967 4951 22973
rect 4893 22933 4905 22967
rect 4939 22964 4951 22967
rect 5442 22964 5448 22976
rect 4939 22936 5448 22964
rect 4939 22933 4951 22936
rect 4893 22927 4951 22933
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 5810 22924 5816 22976
rect 5868 22924 5874 22976
rect 5905 22967 5963 22973
rect 5905 22933 5917 22967
rect 5951 22964 5963 22967
rect 7116 22964 7144 23004
rect 9674 22992 9680 23004
rect 9732 22992 9738 23044
rect 9953 23035 10011 23041
rect 9953 23001 9965 23035
rect 9999 23001 10011 23035
rect 9953 22995 10011 23001
rect 5951 22936 7144 22964
rect 7193 22967 7251 22973
rect 5951 22933 5963 22936
rect 5905 22927 5963 22933
rect 7193 22933 7205 22967
rect 7239 22964 7251 22967
rect 7466 22964 7472 22976
rect 7239 22936 7472 22964
rect 7239 22933 7251 22936
rect 7193 22927 7251 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 8021 22967 8079 22973
rect 8021 22933 8033 22967
rect 8067 22964 8079 22967
rect 8202 22964 8208 22976
rect 8067 22936 8208 22964
rect 8067 22933 8079 22936
rect 8021 22927 8079 22933
rect 8202 22924 8208 22936
rect 8260 22924 8266 22976
rect 9306 22964 9312 22976
rect 9267 22936 9312 22964
rect 9306 22924 9312 22936
rect 9364 22924 9370 22976
rect 9968 22964 9996 22995
rect 10042 22992 10048 23044
rect 10100 23032 10106 23044
rect 10704 23032 10732 23140
rect 11146 23128 11152 23140
rect 11204 23128 11210 23180
rect 11440 23177 11468 23276
rect 14734 23264 14740 23316
rect 14792 23304 14798 23316
rect 15102 23304 15108 23316
rect 14792 23276 15108 23304
rect 14792 23264 14798 23276
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 17678 23264 17684 23316
rect 17736 23304 17742 23316
rect 18325 23307 18383 23313
rect 18325 23304 18337 23307
rect 17736 23276 18337 23304
rect 17736 23264 17742 23276
rect 18325 23273 18337 23276
rect 18371 23273 18383 23307
rect 18325 23267 18383 23273
rect 30469 23307 30527 23313
rect 30469 23273 30481 23307
rect 30515 23304 30527 23307
rect 34514 23304 34520 23316
rect 30515 23276 34520 23304
rect 30515 23273 30527 23276
rect 30469 23267 30527 23273
rect 34514 23264 34520 23276
rect 34572 23264 34578 23316
rect 14366 23236 14372 23248
rect 13096 23208 14372 23236
rect 13096 23177 13124 23208
rect 14366 23196 14372 23208
rect 14424 23196 14430 23248
rect 14826 23196 14832 23248
rect 14884 23236 14890 23248
rect 14884 23208 30696 23236
rect 14884 23196 14890 23208
rect 11425 23171 11483 23177
rect 11425 23137 11437 23171
rect 11471 23137 11483 23171
rect 13081 23171 13139 23177
rect 13081 23168 13093 23171
rect 11425 23131 11483 23137
rect 11900 23140 13093 23168
rect 11241 23035 11299 23041
rect 11241 23032 11253 23035
rect 10100 23004 10145 23032
rect 10704 23004 11253 23032
rect 10100 22992 10106 23004
rect 11241 23001 11253 23004
rect 11287 23001 11299 23035
rect 11241 22995 11299 23001
rect 11900 22964 11928 23140
rect 13081 23137 13093 23140
rect 13127 23137 13139 23171
rect 13081 23131 13139 23137
rect 13262 23128 13268 23180
rect 13320 23168 13326 23180
rect 13320 23140 13768 23168
rect 13320 23128 13326 23140
rect 12526 23100 12532 23112
rect 12487 23072 12532 23100
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 13740 23100 13768 23140
rect 13814 23128 13820 23180
rect 13872 23168 13878 23180
rect 15194 23168 15200 23180
rect 13872 23140 15200 23168
rect 13872 23128 13878 23140
rect 15194 23128 15200 23140
rect 15252 23128 15258 23180
rect 16301 23171 16359 23177
rect 16301 23137 16313 23171
rect 16347 23168 16359 23171
rect 17402 23168 17408 23180
rect 16347 23140 17408 23168
rect 16347 23137 16359 23140
rect 16301 23131 16359 23137
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 19518 23168 19524 23180
rect 19479 23140 19524 23168
rect 19518 23128 19524 23140
rect 19576 23128 19582 23180
rect 18506 23100 18512 23112
rect 13740 23072 14688 23100
rect 18467 23072 18512 23100
rect 13173 23035 13231 23041
rect 13173 23001 13185 23035
rect 13219 23001 13231 23035
rect 13173 22995 13231 23001
rect 13725 23035 13783 23041
rect 13725 23001 13737 23035
rect 13771 23032 13783 23035
rect 14660 23032 14688 23072
rect 18506 23060 18512 23072
rect 18564 23060 18570 23112
rect 23290 23100 23296 23112
rect 23251 23072 23296 23100
rect 23290 23060 23296 23072
rect 23348 23060 23354 23112
rect 30668 23109 30696 23208
rect 30653 23103 30711 23109
rect 30653 23069 30665 23103
rect 30699 23069 30711 23103
rect 30653 23063 30711 23069
rect 15105 23035 15163 23041
rect 15105 23032 15117 23035
rect 13771 23004 14596 23032
rect 14660 23004 15117 23032
rect 13771 23001 13783 23004
rect 13725 22995 13783 23001
rect 9968 22936 11928 22964
rect 12345 22967 12403 22973
rect 12345 22933 12357 22967
rect 12391 22964 12403 22967
rect 12434 22964 12440 22976
rect 12391 22936 12440 22964
rect 12391 22933 12403 22936
rect 12345 22927 12403 22933
rect 12434 22924 12440 22936
rect 12492 22924 12498 22976
rect 13188 22964 13216 22995
rect 14090 22964 14096 22976
rect 13188 22936 14096 22964
rect 14090 22924 14096 22936
rect 14148 22924 14154 22976
rect 14274 22964 14280 22976
rect 14235 22936 14280 22964
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14568 22964 14596 23004
rect 15105 23001 15117 23004
rect 15151 23001 15163 23035
rect 15105 22995 15163 23001
rect 15197 23035 15255 23041
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 15562 23032 15568 23044
rect 15243 23004 15568 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 15562 22992 15568 23004
rect 15620 22992 15626 23044
rect 15749 23035 15807 23041
rect 15749 23001 15761 23035
rect 15795 23001 15807 23035
rect 15749 22995 15807 23001
rect 16393 23035 16451 23041
rect 16393 23001 16405 23035
rect 16439 23032 16451 23035
rect 17126 23032 17132 23044
rect 16439 23004 17132 23032
rect 16439 23001 16451 23004
rect 16393 22995 16451 23001
rect 15654 22964 15660 22976
rect 14568 22936 15660 22964
rect 15654 22924 15660 22936
rect 15712 22924 15718 22976
rect 15764 22964 15792 22995
rect 17126 22992 17132 23004
rect 17184 22992 17190 23044
rect 17310 23032 17316 23044
rect 17271 23004 17316 23032
rect 17310 22992 17316 23004
rect 17368 22992 17374 23044
rect 19613 23035 19671 23041
rect 19613 23001 19625 23035
rect 19659 23001 19671 23035
rect 20162 23032 20168 23044
rect 20123 23004 20168 23032
rect 19613 22995 19671 23001
rect 16758 22964 16764 22976
rect 15764 22936 16764 22964
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 19628 22964 19656 22995
rect 20162 22992 20168 23004
rect 20220 22992 20226 23044
rect 19392 22936 19656 22964
rect 19392 22924 19398 22936
rect 22186 22924 22192 22976
rect 22244 22964 22250 22976
rect 23109 22967 23167 22973
rect 23109 22964 23121 22967
rect 22244 22936 23121 22964
rect 22244 22924 22250 22936
rect 23109 22933 23121 22936
rect 23155 22933 23167 22967
rect 23109 22927 23167 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 3234 22760 3240 22772
rect 1964 22732 3240 22760
rect 1964 22701 1992 22732
rect 3234 22720 3240 22732
rect 3292 22720 3298 22772
rect 4249 22763 4307 22769
rect 4249 22729 4261 22763
rect 4295 22760 4307 22763
rect 8110 22760 8116 22772
rect 4295 22732 8116 22760
rect 4295 22729 4307 22732
rect 4249 22723 4307 22729
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 9950 22760 9956 22772
rect 8404 22732 9956 22760
rect 1949 22695 2007 22701
rect 1949 22661 1961 22695
rect 1995 22661 2007 22695
rect 1949 22655 2007 22661
rect 2774 22652 2780 22704
rect 2832 22692 2838 22704
rect 3053 22695 3111 22701
rect 3053 22692 3065 22695
rect 2832 22664 3065 22692
rect 2832 22652 2838 22664
rect 3053 22661 3065 22664
rect 3099 22661 3111 22695
rect 3053 22655 3111 22661
rect 3145 22695 3203 22701
rect 3145 22661 3157 22695
rect 3191 22692 3203 22695
rect 3510 22692 3516 22704
rect 3191 22664 3516 22692
rect 3191 22661 3203 22664
rect 3145 22655 3203 22661
rect 3510 22652 3516 22664
rect 3568 22652 3574 22704
rect 5169 22695 5227 22701
rect 5169 22661 5181 22695
rect 5215 22692 5227 22695
rect 8404 22692 8432 22732
rect 9950 22720 9956 22732
rect 10008 22720 10014 22772
rect 10042 22720 10048 22772
rect 10100 22760 10106 22772
rect 11793 22763 11851 22769
rect 11793 22760 11805 22763
rect 10100 22732 11805 22760
rect 10100 22720 10106 22732
rect 11793 22729 11805 22732
rect 11839 22729 11851 22763
rect 14274 22760 14280 22772
rect 11793 22723 11851 22729
rect 13740 22732 14280 22760
rect 10134 22692 10140 22704
rect 5215 22664 8432 22692
rect 8496 22664 9904 22692
rect 10095 22664 10140 22692
rect 5215 22661 5227 22664
rect 5169 22655 5227 22661
rect 4157 22627 4215 22633
rect 4157 22593 4169 22627
rect 4203 22593 4215 22627
rect 4157 22587 4215 22593
rect 5077 22627 5135 22633
rect 5077 22593 5089 22627
rect 5123 22624 5135 22627
rect 5534 22624 5540 22636
rect 5123 22596 5540 22624
rect 5123 22593 5135 22596
rect 5077 22587 5135 22593
rect 1857 22559 1915 22565
rect 1857 22525 1869 22559
rect 1903 22525 1915 22559
rect 2130 22556 2136 22568
rect 2091 22528 2136 22556
rect 1857 22519 1915 22525
rect 1872 22488 1900 22519
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 4172 22556 4200 22587
rect 5534 22584 5540 22596
rect 5592 22584 5598 22636
rect 5718 22584 5724 22636
rect 5776 22624 5782 22636
rect 5813 22627 5871 22633
rect 5813 22624 5825 22627
rect 5776 22596 5825 22624
rect 5776 22584 5782 22596
rect 5813 22593 5825 22596
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 5905 22627 5963 22633
rect 5905 22593 5917 22627
rect 5951 22624 5963 22627
rect 5994 22624 6000 22636
rect 5951 22596 6000 22624
rect 5951 22593 5963 22596
rect 5905 22587 5963 22593
rect 5994 22584 6000 22596
rect 6052 22584 6058 22636
rect 6270 22584 6276 22636
rect 6328 22624 6334 22636
rect 6822 22624 6828 22636
rect 6328 22596 6828 22624
rect 6328 22584 6334 22596
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22624 7527 22627
rect 8496 22624 8524 22664
rect 7515 22596 8524 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 8570 22584 8576 22636
rect 8628 22624 8634 22636
rect 8665 22627 8723 22633
rect 8665 22624 8677 22627
rect 8628 22596 8677 22624
rect 8628 22584 8634 22596
rect 8665 22593 8677 22596
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 9122 22584 9128 22636
rect 9180 22624 9186 22636
rect 9309 22627 9367 22633
rect 9309 22624 9321 22627
rect 9180 22596 9321 22624
rect 9180 22584 9186 22596
rect 9309 22593 9321 22596
rect 9355 22593 9367 22627
rect 9309 22587 9367 22593
rect 6086 22556 6092 22568
rect 4172 22528 6092 22556
rect 6086 22516 6092 22528
rect 6144 22516 6150 22568
rect 3605 22491 3663 22497
rect 1872 22460 2912 22488
rect 2884 22429 2912 22460
rect 3605 22457 3617 22491
rect 3651 22488 3663 22491
rect 3786 22488 3792 22500
rect 3651 22460 3792 22488
rect 3651 22457 3663 22460
rect 3605 22451 3663 22457
rect 3786 22448 3792 22460
rect 3844 22488 3850 22500
rect 9876 22488 9904 22664
rect 10134 22652 10140 22664
rect 10192 22652 10198 22704
rect 10226 22652 10232 22704
rect 10284 22692 10290 22704
rect 10686 22692 10692 22704
rect 10284 22664 10692 22692
rect 10284 22652 10290 22664
rect 10686 22652 10692 22664
rect 10744 22652 10750 22704
rect 12618 22692 12624 22704
rect 12579 22664 12624 22692
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 13170 22692 13176 22704
rect 13131 22664 13176 22692
rect 13170 22652 13176 22664
rect 13228 22652 13234 22704
rect 13740 22701 13768 22732
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 15470 22720 15476 22772
rect 15528 22760 15534 22772
rect 29730 22760 29736 22772
rect 15528 22732 29736 22760
rect 15528 22720 15534 22732
rect 29730 22720 29736 22732
rect 29788 22720 29794 22772
rect 13725 22695 13783 22701
rect 13725 22661 13737 22695
rect 13771 22661 13783 22695
rect 13725 22655 13783 22661
rect 13814 22652 13820 22704
rect 13872 22692 13878 22704
rect 13872 22664 13917 22692
rect 13872 22652 13878 22664
rect 14090 22652 14096 22704
rect 14148 22692 14154 22704
rect 16117 22695 16175 22701
rect 16117 22692 16129 22695
rect 14148 22664 16129 22692
rect 14148 22652 14154 22664
rect 16117 22661 16129 22664
rect 16163 22661 16175 22695
rect 16117 22655 16175 22661
rect 11514 22584 11520 22636
rect 11572 22624 11578 22636
rect 11701 22627 11759 22633
rect 11701 22624 11713 22627
rect 11572 22596 11713 22624
rect 11572 22584 11578 22596
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 15381 22627 15439 22633
rect 15381 22593 15393 22627
rect 15427 22593 15439 22627
rect 16022 22624 16028 22636
rect 15983 22596 16028 22624
rect 15381 22587 15439 22593
rect 10045 22559 10103 22565
rect 10045 22525 10057 22559
rect 10091 22556 10103 22559
rect 10778 22556 10784 22568
rect 10091 22528 10784 22556
rect 10091 22525 10103 22528
rect 10045 22519 10103 22525
rect 10778 22516 10784 22528
rect 10836 22516 10842 22568
rect 12529 22559 12587 22565
rect 12529 22525 12541 22559
rect 12575 22556 12587 22559
rect 12710 22556 12716 22568
rect 12575 22528 12716 22556
rect 12575 22525 12587 22528
rect 12529 22519 12587 22525
rect 12710 22516 12716 22528
rect 12768 22516 12774 22568
rect 14366 22556 14372 22568
rect 14327 22528 14372 22556
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 12342 22488 12348 22500
rect 3844 22460 9536 22488
rect 9876 22460 12348 22488
rect 3844 22448 3850 22460
rect 2869 22423 2927 22429
rect 2869 22389 2881 22423
rect 2915 22420 2927 22423
rect 3234 22420 3240 22432
rect 2915 22392 3240 22420
rect 2915 22389 2927 22392
rect 2869 22383 2927 22389
rect 3234 22380 3240 22392
rect 3292 22380 3298 22432
rect 4062 22380 4068 22432
rect 4120 22420 4126 22432
rect 6178 22420 6184 22432
rect 4120 22392 6184 22420
rect 4120 22380 4126 22392
rect 6178 22380 6184 22392
rect 6236 22380 6242 22432
rect 6914 22420 6920 22432
rect 6875 22392 6920 22420
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 7282 22380 7288 22432
rect 7340 22420 7346 22432
rect 7561 22423 7619 22429
rect 7561 22420 7573 22423
rect 7340 22392 7573 22420
rect 7340 22380 7346 22392
rect 7561 22389 7573 22392
rect 7607 22389 7619 22423
rect 8754 22420 8760 22432
rect 8715 22392 8760 22420
rect 7561 22383 7619 22389
rect 8754 22380 8760 22392
rect 8812 22380 8818 22432
rect 9398 22420 9404 22432
rect 9359 22392 9404 22420
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 9508 22420 9536 22460
rect 12342 22448 12348 22460
rect 12400 22448 12406 22500
rect 15396 22488 15424 22587
rect 16022 22584 16028 22596
rect 16080 22584 16086 22636
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22624 18199 22627
rect 21542 22624 21548 22636
rect 18187 22596 21548 22624
rect 18187 22593 18199 22596
rect 18141 22587 18199 22593
rect 21542 22584 21548 22596
rect 21600 22624 21606 22636
rect 23474 22624 23480 22636
rect 21600 22596 23480 22624
rect 21600 22584 21606 22596
rect 23474 22584 23480 22596
rect 23532 22584 23538 22636
rect 36725 22627 36783 22633
rect 36725 22624 36737 22627
rect 31726 22596 36737 22624
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 17586 22556 17592 22568
rect 16632 22528 17592 22556
rect 16632 22516 16638 22528
rect 17586 22516 17592 22528
rect 17644 22556 17650 22568
rect 31726 22556 31754 22596
rect 36725 22593 36737 22596
rect 36771 22593 36783 22627
rect 36725 22587 36783 22593
rect 37826 22584 37832 22636
rect 37884 22624 37890 22636
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 37884 22596 38025 22624
rect 37884 22584 37890 22596
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 17644 22528 31754 22556
rect 17644 22516 17650 22528
rect 38194 22488 38200 22500
rect 13188 22460 15424 22488
rect 38155 22460 38200 22488
rect 9858 22420 9864 22432
rect 9508 22392 9864 22420
rect 9858 22380 9864 22392
rect 9916 22380 9922 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10502 22420 10508 22432
rect 10008 22392 10508 22420
rect 10008 22380 10014 22392
rect 10502 22380 10508 22392
rect 10560 22380 10566 22432
rect 12894 22380 12900 22432
rect 12952 22420 12958 22432
rect 13188 22420 13216 22460
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 12952 22392 13216 22420
rect 12952 22380 12958 22392
rect 15194 22380 15200 22432
rect 15252 22420 15258 22432
rect 15473 22423 15531 22429
rect 15473 22420 15485 22423
rect 15252 22392 15485 22420
rect 15252 22380 15258 22392
rect 15473 22389 15485 22392
rect 15519 22389 15531 22423
rect 15473 22383 15531 22389
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 18233 22423 18291 22429
rect 18233 22420 18245 22423
rect 18012 22392 18245 22420
rect 18012 22380 18018 22392
rect 18233 22389 18245 22392
rect 18279 22389 18291 22423
rect 18233 22383 18291 22389
rect 36817 22423 36875 22429
rect 36817 22389 36829 22423
rect 36863 22420 36875 22423
rect 38010 22420 38016 22432
rect 36863 22392 38016 22420
rect 36863 22389 36875 22392
rect 36817 22383 36875 22389
rect 38010 22380 38016 22392
rect 38068 22380 38074 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3234 22176 3240 22228
rect 3292 22216 3298 22228
rect 3292 22188 9674 22216
rect 3292 22176 3298 22188
rect 2498 22108 2504 22160
rect 2556 22148 2562 22160
rect 4798 22148 4804 22160
rect 2556 22120 4804 22148
rect 2556 22108 2562 22120
rect 4798 22108 4804 22120
rect 4856 22108 4862 22160
rect 8386 22108 8392 22160
rect 8444 22148 8450 22160
rect 8481 22151 8539 22157
rect 8481 22148 8493 22151
rect 8444 22120 8493 22148
rect 8444 22108 8450 22120
rect 8481 22117 8493 22120
rect 8527 22117 8539 22151
rect 9646 22148 9674 22188
rect 9858 22176 9864 22228
rect 9916 22216 9922 22228
rect 15010 22216 15016 22228
rect 9916 22188 15016 22216
rect 9916 22176 9922 22188
rect 15010 22176 15016 22188
rect 15068 22176 15074 22228
rect 15378 22176 15384 22228
rect 15436 22216 15442 22228
rect 15746 22216 15752 22228
rect 15436 22188 15752 22216
rect 15436 22176 15442 22188
rect 15746 22176 15752 22188
rect 15804 22176 15810 22228
rect 20254 22216 20260 22228
rect 19996 22188 20260 22216
rect 15286 22148 15292 22160
rect 9646 22120 15292 22148
rect 8481 22111 8539 22117
rect 15286 22108 15292 22120
rect 15344 22108 15350 22160
rect 16758 22108 16764 22160
rect 16816 22148 16822 22160
rect 18785 22151 18843 22157
rect 18785 22148 18797 22151
rect 16816 22120 18797 22148
rect 16816 22108 16822 22120
rect 3234 22040 3240 22092
rect 3292 22080 3298 22092
rect 3602 22080 3608 22092
rect 3292 22052 3608 22080
rect 3292 22040 3298 22052
rect 3602 22040 3608 22052
rect 3660 22040 3666 22092
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 4632 22052 6285 22080
rect 4632 22024 4660 22052
rect 6273 22049 6285 22052
rect 6319 22049 6331 22083
rect 9140 22080 9444 22092
rect 10042 22080 10048 22092
rect 6273 22043 6331 22049
rect 9048 22064 10048 22080
rect 9048 22052 9168 22064
rect 9416 22052 10048 22064
rect 1578 22012 1584 22024
rect 1539 21984 1584 22012
rect 1578 21972 1584 21984
rect 1636 21972 1642 22024
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 3970 22012 3976 22024
rect 1903 21984 3976 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 3970 21972 3976 21984
rect 4028 21972 4034 22024
rect 4246 22012 4252 22024
rect 4207 21984 4252 22012
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 4614 21972 4620 22024
rect 4672 21972 4678 22024
rect 4893 22015 4951 22021
rect 4893 21981 4905 22015
rect 4939 22012 4951 22015
rect 5074 22012 5080 22024
rect 4939 21984 5080 22012
rect 4939 21981 4951 21984
rect 4893 21975 4951 21981
rect 5074 21972 5080 21984
rect 5132 21972 5138 22024
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 22012 5595 22015
rect 6181 22015 6239 22021
rect 5583 21984 6132 22012
rect 5583 21981 5595 21984
rect 5537 21975 5595 21981
rect 2958 21944 2964 21956
rect 2919 21916 2964 21944
rect 2958 21904 2964 21916
rect 3016 21904 3022 21956
rect 4341 21947 4399 21953
rect 4341 21913 4353 21947
rect 4387 21944 4399 21947
rect 4430 21944 4436 21956
rect 4387 21916 4436 21944
rect 4387 21913 4399 21916
rect 4341 21907 4399 21913
rect 4430 21904 4436 21916
rect 4488 21904 4494 21956
rect 5718 21944 5724 21956
rect 5552 21916 5724 21944
rect 3053 21879 3111 21885
rect 3053 21845 3065 21879
rect 3099 21876 3111 21879
rect 3234 21876 3240 21888
rect 3099 21848 3240 21876
rect 3099 21845 3111 21848
rect 3053 21839 3111 21845
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4706 21876 4712 21888
rect 4212 21848 4712 21876
rect 4212 21836 4218 21848
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 4985 21879 5043 21885
rect 4985 21845 4997 21879
rect 5031 21876 5043 21879
rect 5552 21876 5580 21916
rect 5718 21904 5724 21916
rect 5776 21904 5782 21956
rect 5031 21848 5580 21876
rect 5629 21879 5687 21885
rect 5031 21845 5043 21848
rect 4985 21839 5043 21845
rect 5629 21845 5641 21879
rect 5675 21876 5687 21879
rect 5902 21876 5908 21888
rect 5675 21848 5908 21876
rect 5675 21845 5687 21848
rect 5629 21839 5687 21845
rect 5902 21836 5908 21848
rect 5960 21836 5966 21888
rect 6104 21876 6132 21984
rect 6181 21981 6193 22015
rect 6227 22012 6239 22015
rect 6546 22012 6552 22024
rect 6227 21984 6552 22012
rect 6227 21981 6239 21984
rect 6181 21975 6239 21981
rect 6546 21972 6552 21984
rect 6604 21972 6610 22024
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 7650 22012 7656 22024
rect 7101 21975 7159 21981
rect 7208 21984 7656 22012
rect 7006 21904 7012 21956
rect 7064 21944 7070 21956
rect 7116 21944 7144 21975
rect 7208 21953 7236 21984
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 22012 7803 22015
rect 8110 22012 8116 22024
rect 7791 21984 8116 22012
rect 7791 21981 7803 21984
rect 7745 21975 7803 21981
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 8413 22015 8471 22021
rect 8413 21981 8425 22015
rect 8459 22012 8471 22015
rect 9048 22012 9076 22052
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 10229 22083 10287 22089
rect 10229 22049 10241 22083
rect 10275 22080 10287 22083
rect 11790 22080 11796 22092
rect 10275 22052 11796 22080
rect 10275 22049 10287 22052
rect 10229 22043 10287 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 11882 22040 11888 22092
rect 11940 22080 11946 22092
rect 15102 22080 15108 22092
rect 11940 22052 14320 22080
rect 15063 22052 15108 22080
rect 11940 22040 11946 22052
rect 8459 21984 9076 22012
rect 8459 21981 8471 21984
rect 8413 21975 8471 21981
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12894 22012 12900 22024
rect 12492 21984 12537 22012
rect 12855 21984 12900 22012
rect 12492 21972 12498 21984
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 13262 21972 13268 22024
rect 13320 22012 13326 22024
rect 13320 21988 13492 22012
rect 13549 22009 13607 22015
rect 13549 21988 13561 22009
rect 13320 21984 13561 21988
rect 13320 21972 13326 21984
rect 13464 21975 13561 21984
rect 13595 21975 13607 22009
rect 14292 22014 14320 22052
rect 15102 22040 15108 22052
rect 15160 22040 15166 22092
rect 15930 22080 15936 22092
rect 15891 22052 15936 22080
rect 15930 22040 15936 22052
rect 15988 22040 15994 22092
rect 17034 22080 17040 22092
rect 16995 22052 17040 22080
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 17328 22089 17356 22120
rect 18785 22117 18797 22120
rect 18831 22117 18843 22151
rect 18785 22111 18843 22117
rect 17313 22083 17371 22089
rect 17313 22049 17325 22083
rect 17359 22080 17371 22083
rect 18233 22083 18291 22089
rect 17359 22052 17393 22080
rect 17359 22049 17371 22052
rect 17313 22043 17371 22049
rect 18233 22049 18245 22083
rect 18279 22080 18291 22083
rect 19996 22080 20024 22188
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 37826 22216 37832 22228
rect 37787 22188 37832 22216
rect 37826 22176 37832 22188
rect 37884 22176 37890 22228
rect 20162 22108 20168 22160
rect 20220 22148 20226 22160
rect 20346 22148 20352 22160
rect 20220 22120 20352 22148
rect 20220 22108 20226 22120
rect 20346 22108 20352 22120
rect 20404 22148 20410 22160
rect 20625 22151 20683 22157
rect 20625 22148 20637 22151
rect 20404 22120 20637 22148
rect 20404 22108 20410 22120
rect 20625 22117 20637 22120
rect 20671 22117 20683 22151
rect 20625 22111 20683 22117
rect 18279 22052 20024 22080
rect 20073 22083 20131 22089
rect 18279 22049 18291 22052
rect 18233 22043 18291 22049
rect 20073 22049 20085 22083
rect 20119 22080 20131 22083
rect 23106 22080 23112 22092
rect 20119 22052 23112 22080
rect 20119 22049 20131 22052
rect 20073 22043 20131 22049
rect 23106 22040 23112 22052
rect 23164 22040 23170 22092
rect 25317 22083 25375 22089
rect 25317 22049 25329 22083
rect 25363 22080 25375 22083
rect 28994 22080 29000 22092
rect 25363 22052 29000 22080
rect 25363 22049 25375 22052
rect 25317 22043 25375 22049
rect 28994 22040 29000 22052
rect 29052 22040 29058 22092
rect 14369 22015 14427 22021
rect 14369 22014 14381 22015
rect 14292 21986 14381 22014
rect 14369 21981 14381 21986
rect 14415 21981 14427 22015
rect 38010 22012 38016 22024
rect 37971 21984 38016 22012
rect 14369 21975 14427 21981
rect 13464 21969 13607 21975
rect 38010 21972 38016 21984
rect 38068 21972 38074 22024
rect 13464 21960 13584 21969
rect 7064 21916 7144 21944
rect 7193 21947 7251 21953
rect 7064 21904 7070 21916
rect 7193 21913 7205 21947
rect 7239 21913 7251 21947
rect 9214 21944 9220 21956
rect 9175 21916 9220 21944
rect 7193 21907 7251 21913
rect 9214 21904 9220 21916
rect 9272 21904 9278 21956
rect 9306 21904 9312 21956
rect 9364 21944 9370 21956
rect 10778 21944 10784 21956
rect 9364 21916 9409 21944
rect 10739 21916 10784 21944
rect 9364 21904 9370 21916
rect 10778 21904 10784 21916
rect 10836 21904 10842 21956
rect 10870 21904 10876 21956
rect 10928 21944 10934 21956
rect 11422 21944 11428 21956
rect 10928 21916 10973 21944
rect 11383 21916 11428 21944
rect 10928 21904 10934 21916
rect 11422 21904 11428 21916
rect 11480 21904 11486 21956
rect 13633 21947 13691 21953
rect 13633 21913 13645 21947
rect 13679 21944 13691 21947
rect 14550 21944 14556 21956
rect 13679 21916 14556 21944
rect 13679 21913 13691 21916
rect 13633 21907 13691 21913
rect 14550 21904 14556 21916
rect 14608 21904 14614 21956
rect 15194 21904 15200 21956
rect 15252 21944 15258 21956
rect 17129 21947 17187 21953
rect 15252 21916 15297 21944
rect 15252 21904 15258 21916
rect 17129 21913 17141 21947
rect 17175 21913 17187 21947
rect 17129 21907 17187 21913
rect 18325 21947 18383 21953
rect 18325 21913 18337 21947
rect 18371 21944 18383 21947
rect 19150 21944 19156 21956
rect 18371 21916 19156 21944
rect 18371 21913 18383 21916
rect 18325 21907 18383 21913
rect 6546 21876 6552 21888
rect 6104 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 7558 21836 7564 21888
rect 7616 21876 7622 21888
rect 7837 21879 7895 21885
rect 7837 21876 7849 21879
rect 7616 21848 7849 21876
rect 7616 21836 7622 21848
rect 7837 21845 7849 21848
rect 7883 21845 7895 21879
rect 7837 21839 7895 21845
rect 8294 21836 8300 21888
rect 8352 21876 8358 21888
rect 11882 21876 11888 21888
rect 8352 21848 11888 21876
rect 8352 21836 8358 21848
rect 11882 21836 11888 21848
rect 11940 21836 11946 21888
rect 12250 21876 12256 21888
rect 12211 21848 12256 21876
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 12989 21879 13047 21885
rect 12989 21845 13001 21879
rect 13035 21876 13047 21879
rect 14274 21876 14280 21888
rect 13035 21848 14280 21876
rect 13035 21845 13047 21848
rect 12989 21839 13047 21845
rect 14274 21836 14280 21848
rect 14332 21836 14338 21888
rect 14458 21876 14464 21888
rect 14419 21848 14464 21876
rect 14458 21836 14464 21848
rect 14516 21836 14522 21888
rect 17144 21876 17172 21907
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 20165 21947 20223 21953
rect 20165 21913 20177 21947
rect 20211 21944 20223 21947
rect 20530 21944 20536 21956
rect 20211 21916 20536 21944
rect 20211 21913 20223 21916
rect 20165 21907 20223 21913
rect 20530 21904 20536 21916
rect 20588 21904 20594 21956
rect 25406 21904 25412 21956
rect 25464 21944 25470 21956
rect 26329 21947 26387 21953
rect 26329 21944 26341 21947
rect 25464 21916 25509 21944
rect 26160 21916 26341 21944
rect 25464 21904 25470 21916
rect 19426 21876 19432 21888
rect 17144 21848 19432 21876
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 21726 21876 21732 21888
rect 21687 21848 21732 21876
rect 21726 21836 21732 21848
rect 21784 21836 21790 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 26160 21876 26188 21916
rect 26329 21913 26341 21916
rect 26375 21913 26387 21947
rect 26329 21907 26387 21913
rect 22612 21848 26188 21876
rect 22612 21836 22618 21848
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 3234 21632 3240 21684
rect 3292 21672 3298 21684
rect 3970 21672 3976 21684
rect 3292 21644 3976 21672
rect 3292 21632 3298 21644
rect 3970 21632 3976 21644
rect 4028 21632 4034 21684
rect 4890 21672 4896 21684
rect 4724 21644 4896 21672
rect 1854 21604 1860 21616
rect 1815 21576 1860 21604
rect 1854 21564 1860 21576
rect 1912 21564 1918 21616
rect 3421 21607 3479 21613
rect 3421 21573 3433 21607
rect 3467 21604 3479 21607
rect 4154 21604 4160 21616
rect 3467 21576 4160 21604
rect 3467 21573 3479 21576
rect 3421 21567 3479 21573
rect 4154 21564 4160 21576
rect 4212 21564 4218 21616
rect 4617 21607 4675 21613
rect 4617 21573 4629 21607
rect 4663 21604 4675 21607
rect 4724 21604 4752 21644
rect 4890 21632 4896 21644
rect 4948 21632 4954 21684
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5905 21675 5963 21681
rect 5905 21672 5917 21675
rect 5132 21644 5917 21672
rect 5132 21632 5138 21644
rect 5905 21641 5917 21644
rect 5951 21641 5963 21675
rect 11054 21672 11060 21684
rect 5905 21635 5963 21641
rect 8036 21644 11060 21672
rect 7190 21604 7196 21616
rect 4663 21576 4752 21604
rect 7151 21576 7196 21604
rect 4663 21573 4675 21576
rect 4617 21567 4675 21573
rect 7190 21564 7196 21576
rect 7248 21564 7254 21616
rect 7285 21607 7343 21613
rect 7285 21573 7297 21607
rect 7331 21604 7343 21607
rect 7374 21604 7380 21616
rect 7331 21576 7380 21604
rect 7331 21573 7343 21576
rect 7285 21567 7343 21573
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 5813 21539 5871 21545
rect 4172 21508 4384 21536
rect 1765 21471 1823 21477
rect 1765 21437 1777 21471
rect 1811 21468 1823 21471
rect 2777 21471 2835 21477
rect 1811 21440 2728 21468
rect 1811 21437 1823 21440
rect 1765 21431 1823 21437
rect 2700 21332 2728 21440
rect 2777 21437 2789 21471
rect 2823 21437 2835 21471
rect 2777 21431 2835 21437
rect 3329 21471 3387 21477
rect 3329 21437 3341 21471
rect 3375 21468 3387 21471
rect 3602 21468 3608 21480
rect 3375 21440 3608 21468
rect 3375 21437 3387 21440
rect 3329 21431 3387 21437
rect 2792 21400 2820 21431
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 3786 21468 3792 21480
rect 3747 21440 3792 21468
rect 3786 21428 3792 21440
rect 3844 21428 3850 21480
rect 4172 21400 4200 21508
rect 4356 21468 4384 21508
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 6822 21536 6828 21548
rect 5859 21508 6828 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 6822 21496 6828 21508
rect 6880 21496 6886 21548
rect 4525 21471 4583 21477
rect 4525 21468 4537 21471
rect 4356 21440 4537 21468
rect 4525 21437 4537 21440
rect 4571 21468 4583 21471
rect 7469 21471 7527 21477
rect 7469 21468 7481 21471
rect 4571 21440 7481 21468
rect 4571 21437 4583 21440
rect 4525 21431 4583 21437
rect 7469 21437 7481 21440
rect 7515 21468 7527 21471
rect 8036 21468 8064 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11422 21632 11428 21684
rect 11480 21672 11486 21684
rect 25225 21675 25283 21681
rect 11480 21644 22048 21672
rect 11480 21632 11486 21644
rect 8849 21607 8907 21613
rect 8849 21573 8861 21607
rect 8895 21604 8907 21607
rect 9766 21604 9772 21616
rect 8895 21576 9772 21604
rect 8895 21573 8907 21576
rect 8849 21567 8907 21573
rect 9766 21564 9772 21576
rect 9824 21564 9830 21616
rect 9858 21564 9864 21616
rect 9916 21604 9922 21616
rect 11606 21604 11612 21616
rect 9916 21576 11612 21604
rect 9916 21564 9922 21576
rect 11606 21564 11612 21576
rect 11664 21564 11670 21616
rect 12161 21607 12219 21613
rect 12161 21573 12173 21607
rect 12207 21604 12219 21607
rect 12250 21604 12256 21616
rect 12207 21576 12256 21604
rect 12207 21573 12219 21576
rect 12161 21567 12219 21573
rect 12250 21564 12256 21576
rect 12308 21564 12314 21616
rect 13357 21607 13415 21613
rect 13357 21573 13369 21607
rect 13403 21604 13415 21607
rect 14458 21604 14464 21616
rect 13403 21576 14464 21604
rect 13403 21573 13415 21576
rect 13357 21567 13415 21573
rect 14458 21564 14464 21576
rect 14516 21564 14522 21616
rect 17126 21564 17132 21616
rect 17184 21604 17190 21616
rect 18509 21607 18567 21613
rect 18509 21604 18521 21607
rect 17184 21576 18521 21604
rect 17184 21564 17190 21576
rect 18509 21573 18521 21576
rect 18555 21573 18567 21607
rect 19150 21604 19156 21616
rect 19111 21576 19156 21604
rect 18509 21567 18567 21573
rect 19150 21564 19156 21576
rect 19208 21564 19214 21616
rect 19889 21607 19947 21613
rect 19889 21573 19901 21607
rect 19935 21604 19947 21607
rect 19978 21604 19984 21616
rect 19935 21576 19984 21604
rect 19935 21573 19947 21576
rect 19889 21567 19947 21573
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 22020 21604 22048 21644
rect 25225 21641 25237 21675
rect 25271 21672 25283 21675
rect 25406 21672 25412 21684
rect 25271 21644 25412 21672
rect 25271 21641 25283 21644
rect 25225 21635 25283 21641
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 32306 21672 32312 21684
rect 32267 21644 32312 21672
rect 32306 21632 32312 21644
rect 32364 21632 32370 21684
rect 25961 21607 26019 21613
rect 25961 21604 25973 21607
rect 22020 21576 25973 21604
rect 25961 21573 25973 21576
rect 26007 21573 26019 21607
rect 25961 21567 26019 21573
rect 26053 21607 26111 21613
rect 26053 21573 26065 21607
rect 26099 21604 26111 21607
rect 26234 21604 26240 21616
rect 26099 21576 26240 21604
rect 26099 21573 26111 21576
rect 26053 21567 26111 21573
rect 26234 21564 26240 21576
rect 26292 21564 26298 21616
rect 10321 21539 10379 21545
rect 10321 21505 10333 21539
rect 10367 21505 10379 21539
rect 10321 21499 10379 21505
rect 7515 21440 8064 21468
rect 8757 21471 8815 21477
rect 7515 21437 7527 21440
rect 7469 21431 7527 21437
rect 8757 21437 8769 21471
rect 8803 21468 8815 21471
rect 8846 21468 8852 21480
rect 8803 21440 8852 21468
rect 8803 21437 8815 21440
rect 8757 21431 8815 21437
rect 8846 21428 8852 21440
rect 8904 21428 8910 21480
rect 8938 21428 8944 21480
rect 8996 21468 9002 21480
rect 9033 21471 9091 21477
rect 9033 21468 9045 21471
rect 8996 21440 9045 21468
rect 8996 21428 9002 21440
rect 9033 21437 9045 21440
rect 9079 21437 9091 21471
rect 10336 21468 10364 21499
rect 10594 21496 10600 21548
rect 10652 21536 10658 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 10652 21508 10977 21536
rect 10652 21496 10658 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14369 21539 14427 21545
rect 14369 21536 14381 21539
rect 14240 21508 14381 21536
rect 14240 21496 14246 21508
rect 14369 21505 14381 21508
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 14918 21496 14924 21548
rect 14976 21536 14982 21548
rect 15933 21539 15991 21545
rect 15933 21536 15945 21539
rect 14976 21508 15945 21536
rect 14976 21496 14982 21508
rect 15933 21505 15945 21508
rect 15979 21505 15991 21539
rect 15933 21499 15991 21505
rect 18417 21539 18475 21545
rect 18417 21505 18429 21539
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 9033 21431 9091 21437
rect 9140 21440 10364 21468
rect 2792 21372 4200 21400
rect 4706 21360 4712 21412
rect 4764 21400 4770 21412
rect 5077 21403 5135 21409
rect 5077 21400 5089 21403
rect 4764 21372 5089 21400
rect 4764 21360 4770 21372
rect 5077 21369 5089 21372
rect 5123 21369 5135 21403
rect 5077 21363 5135 21369
rect 7282 21360 7288 21412
rect 7340 21400 7346 21412
rect 9140 21400 9168 21440
rect 11146 21428 11152 21480
rect 11204 21468 11210 21480
rect 11882 21468 11888 21480
rect 11204 21440 11888 21468
rect 11204 21428 11210 21440
rect 11882 21428 11888 21440
rect 11940 21428 11946 21480
rect 12069 21471 12127 21477
rect 12069 21437 12081 21471
rect 12115 21468 12127 21471
rect 12710 21468 12716 21480
rect 12115 21440 12716 21468
rect 12115 21437 12127 21440
rect 12069 21431 12127 21437
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 13262 21468 13268 21480
rect 13223 21440 13268 21468
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 16114 21468 16120 21480
rect 14599 21440 16120 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 18432 21468 18460 21499
rect 18598 21496 18604 21548
rect 18656 21536 18662 21548
rect 19061 21539 19119 21545
rect 19061 21536 19073 21539
rect 18656 21508 19073 21536
rect 18656 21496 18662 21508
rect 19061 21505 19073 21508
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21784 21508 22017 21536
rect 21784 21496 21790 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22186 21536 22192 21548
rect 22147 21508 22192 21536
rect 22005 21499 22063 21505
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 23382 21536 23388 21548
rect 23032 21508 23388 21536
rect 19794 21468 19800 21480
rect 18380 21440 18460 21468
rect 19755 21440 19800 21468
rect 18380 21428 18386 21440
rect 19794 21428 19800 21440
rect 19852 21428 19858 21480
rect 7340 21372 9168 21400
rect 7340 21360 7346 21372
rect 9306 21360 9312 21412
rect 9364 21400 9370 21412
rect 12621 21403 12679 21409
rect 9364 21372 12434 21400
rect 9364 21360 9370 21372
rect 4522 21332 4528 21344
rect 2700 21304 4528 21332
rect 4522 21292 4528 21304
rect 4580 21292 4586 21344
rect 6270 21292 6276 21344
rect 6328 21332 6334 21344
rect 9490 21332 9496 21344
rect 6328 21304 9496 21332
rect 6328 21292 6334 21304
rect 9490 21292 9496 21304
rect 9548 21292 9554 21344
rect 10413 21335 10471 21341
rect 10413 21301 10425 21335
rect 10459 21332 10471 21335
rect 10870 21332 10876 21344
rect 10459 21304 10876 21332
rect 10459 21301 10471 21304
rect 10413 21295 10471 21301
rect 10870 21292 10876 21304
rect 10928 21292 10934 21344
rect 11057 21335 11115 21341
rect 11057 21301 11069 21335
rect 11103 21332 11115 21335
rect 12158 21332 12164 21344
rect 11103 21304 12164 21332
rect 11103 21301 11115 21304
rect 11057 21295 11115 21301
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 12406 21332 12434 21372
rect 12621 21369 12633 21403
rect 12667 21400 12679 21403
rect 12986 21400 12992 21412
rect 12667 21372 12992 21400
rect 12667 21369 12679 21372
rect 12621 21363 12679 21369
rect 12986 21360 12992 21372
rect 13044 21360 13050 21412
rect 13630 21360 13636 21412
rect 13688 21400 13694 21412
rect 13817 21403 13875 21409
rect 13817 21400 13829 21403
rect 13688 21372 13829 21400
rect 13688 21360 13694 21372
rect 13817 21369 13829 21372
rect 13863 21369 13875 21403
rect 13817 21363 13875 21369
rect 15013 21403 15071 21409
rect 15013 21369 15025 21403
rect 15059 21400 15071 21403
rect 15059 21372 19334 21400
rect 15059 21369 15071 21372
rect 15013 21363 15071 21369
rect 14366 21332 14372 21344
rect 12406 21304 14372 21332
rect 14366 21292 14372 21304
rect 14424 21292 14430 21344
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 16025 21335 16083 21341
rect 16025 21332 16037 21335
rect 15528 21304 16037 21332
rect 15528 21292 15534 21304
rect 16025 21301 16037 21304
rect 16071 21301 16083 21335
rect 16025 21295 16083 21301
rect 16850 21292 16856 21344
rect 16908 21332 16914 21344
rect 18598 21332 18604 21344
rect 16908 21304 18604 21332
rect 16908 21292 16914 21304
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 19306 21332 19334 21372
rect 20346 21360 20352 21412
rect 20404 21400 20410 21412
rect 23032 21400 23060 21508
rect 23382 21496 23388 21508
rect 23440 21536 23446 21548
rect 23753 21539 23811 21545
rect 23753 21536 23765 21539
rect 23440 21508 23765 21536
rect 23440 21496 23446 21508
rect 23753 21505 23765 21508
rect 23799 21505 23811 21539
rect 25130 21536 25136 21548
rect 25091 21508 25136 21536
rect 23753 21499 23811 21505
rect 25130 21496 25136 21508
rect 25188 21496 25194 21548
rect 30466 21496 30472 21548
rect 30524 21536 30530 21548
rect 32493 21539 32551 21545
rect 32493 21536 32505 21539
rect 30524 21508 32505 21536
rect 30524 21496 30530 21508
rect 32493 21505 32505 21508
rect 32539 21505 32551 21539
rect 38010 21536 38016 21548
rect 37971 21508 38016 21536
rect 32493 21499 32551 21505
rect 38010 21496 38016 21508
rect 38068 21496 38074 21548
rect 23106 21428 23112 21480
rect 23164 21468 23170 21480
rect 23293 21471 23351 21477
rect 23164 21440 23257 21468
rect 23164 21428 23170 21440
rect 23293 21437 23305 21471
rect 23339 21468 23351 21471
rect 23658 21468 23664 21480
rect 23339 21440 23664 21468
rect 23339 21437 23351 21440
rect 23293 21431 23351 21437
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 20404 21372 20449 21400
rect 22204 21372 23060 21400
rect 20404 21360 20410 21372
rect 22204 21332 22232 21372
rect 22370 21332 22376 21344
rect 19306 21304 22232 21332
rect 22331 21304 22376 21332
rect 22370 21292 22376 21304
rect 22428 21292 22434 21344
rect 23124 21332 23152 21428
rect 26326 21400 26332 21412
rect 23860 21372 26332 21400
rect 23860 21332 23888 21372
rect 26326 21360 26332 21372
rect 26384 21360 26390 21412
rect 26510 21400 26516 21412
rect 26471 21372 26516 21400
rect 26510 21360 26516 21372
rect 26568 21360 26574 21412
rect 32398 21400 32404 21412
rect 31726 21372 32404 21400
rect 23124 21304 23888 21332
rect 24394 21292 24400 21344
rect 24452 21332 24458 21344
rect 31726 21332 31754 21372
rect 32398 21360 32404 21372
rect 32456 21360 32462 21412
rect 38194 21332 38200 21344
rect 24452 21304 31754 21332
rect 38155 21304 38200 21332
rect 24452 21292 24458 21304
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1854 21088 1860 21140
rect 1912 21128 1918 21140
rect 2130 21128 2136 21140
rect 1912 21100 2136 21128
rect 1912 21088 1918 21100
rect 2130 21088 2136 21100
rect 2188 21128 2194 21140
rect 2188 21100 2912 21128
rect 2188 21088 2194 21100
rect 2774 21060 2780 21072
rect 2746 21020 2780 21060
rect 2832 21020 2838 21072
rect 2884 21060 2912 21100
rect 3234 21088 3240 21140
rect 3292 21128 3298 21140
rect 3292 21100 7604 21128
rect 3292 21088 3298 21100
rect 4706 21060 4712 21072
rect 2884 21032 4712 21060
rect 2225 20995 2283 21001
rect 2225 20961 2237 20995
rect 2271 20992 2283 20995
rect 2746 20992 2774 21020
rect 2884 21001 2912 21032
rect 4706 21020 4712 21032
rect 4764 21020 4770 21072
rect 5261 21063 5319 21069
rect 5261 21029 5273 21063
rect 5307 21060 5319 21063
rect 7466 21060 7472 21072
rect 5307 21032 7472 21060
rect 5307 21029 5319 21032
rect 5261 21023 5319 21029
rect 7466 21020 7472 21032
rect 7524 21020 7530 21072
rect 7576 21060 7604 21100
rect 8938 21088 8944 21140
rect 8996 21128 9002 21140
rect 9306 21128 9312 21140
rect 8996 21100 9312 21128
rect 8996 21088 9002 21100
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 9401 21131 9459 21137
rect 9401 21097 9413 21131
rect 9447 21128 9459 21131
rect 9582 21128 9588 21140
rect 9447 21100 9588 21128
rect 9447 21097 9459 21100
rect 9401 21091 9459 21097
rect 9582 21088 9588 21100
rect 9640 21088 9646 21140
rect 11514 21088 11520 21140
rect 11572 21128 11578 21140
rect 16114 21128 16120 21140
rect 11572 21100 15976 21128
rect 16075 21100 16120 21128
rect 11572 21088 11578 21100
rect 9950 21060 9956 21072
rect 7576 21032 9956 21060
rect 9950 21020 9956 21032
rect 10008 21020 10014 21072
rect 11330 21060 11336 21072
rect 10060 21032 11336 21060
rect 2271 20964 2774 20992
rect 2869 20995 2927 21001
rect 2271 20961 2283 20964
rect 2225 20955 2283 20961
rect 2869 20961 2881 20995
rect 2915 20961 2927 20995
rect 6178 20992 6184 21004
rect 2869 20955 2927 20961
rect 3988 20964 6184 20992
rect 3988 20933 4016 20964
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6549 20995 6607 21001
rect 6549 20961 6561 20995
rect 6595 20992 6607 20995
rect 8662 20992 8668 21004
rect 6595 20964 8668 20992
rect 6595 20961 6607 20964
rect 6549 20955 6607 20961
rect 8662 20952 8668 20964
rect 8720 20952 8726 21004
rect 9766 20992 9772 21004
rect 9048 20964 9772 20992
rect 3973 20927 4031 20933
rect 3973 20893 3985 20927
rect 4019 20893 4031 20927
rect 3973 20887 4031 20893
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 9048 20924 9076 20964
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 10060 21001 10088 21032
rect 11330 21020 11336 21032
rect 11388 21020 11394 21072
rect 12618 21020 12624 21072
rect 12676 21060 12682 21072
rect 12894 21060 12900 21072
rect 12676 21032 12900 21060
rect 12676 21020 12682 21032
rect 12894 21020 12900 21032
rect 12952 21020 12958 21072
rect 13262 21020 13268 21072
rect 13320 21060 13326 21072
rect 14090 21060 14096 21072
rect 13320 21032 14096 21060
rect 13320 21020 13326 21032
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 14366 21020 14372 21072
rect 14424 21060 14430 21072
rect 15838 21060 15844 21072
rect 14424 21032 15844 21060
rect 14424 21020 14430 21032
rect 15838 21020 15844 21032
rect 15896 21020 15902 21072
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20961 10103 20995
rect 10962 20992 10968 21004
rect 10923 20964 10968 20992
rect 10045 20955 10103 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 12529 20995 12587 21001
rect 12529 20961 12541 20995
rect 12575 20992 12587 20995
rect 13170 20992 13176 21004
rect 12575 20964 13176 20992
rect 12575 20961 12587 20964
rect 12529 20955 12587 20961
rect 13170 20952 13176 20964
rect 13228 20992 13234 21004
rect 13630 20992 13636 21004
rect 13228 20964 13636 20992
rect 13228 20952 13234 20964
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 14642 20992 14648 21004
rect 14603 20964 14648 20992
rect 14642 20952 14648 20964
rect 14700 20992 14706 21004
rect 15010 20992 15016 21004
rect 14700 20964 15016 20992
rect 14700 20952 14706 20964
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 15948 20992 15976 21100
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 16206 21088 16212 21140
rect 16264 21128 16270 21140
rect 20530 21128 20536 21140
rect 16264 21100 17908 21128
rect 20491 21100 20536 21128
rect 16264 21088 16270 21100
rect 16022 21020 16028 21072
rect 16080 21060 16086 21072
rect 17880 21060 17908 21100
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 26234 21128 26240 21140
rect 22066 21100 24256 21128
rect 26195 21100 26240 21128
rect 22066 21060 22094 21100
rect 16080 21032 17540 21060
rect 17880 21032 22094 21060
rect 16080 21020 16086 21032
rect 16942 20992 16948 21004
rect 15120 20964 15792 20992
rect 15948 20964 16948 20992
rect 8444 20896 9076 20924
rect 9309 20927 9367 20933
rect 8444 20884 8450 20896
rect 9309 20893 9321 20927
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 2314 20816 2320 20868
rect 2372 20856 2378 20868
rect 2372 20828 2417 20856
rect 2372 20816 2378 20828
rect 4522 20816 4528 20868
rect 4580 20856 4586 20868
rect 4709 20859 4767 20865
rect 4709 20856 4721 20859
rect 4580 20828 4721 20856
rect 4580 20816 4586 20828
rect 4709 20825 4721 20828
rect 4755 20825 4767 20859
rect 4709 20819 4767 20825
rect 4798 20816 4804 20868
rect 4856 20856 4862 20868
rect 5902 20856 5908 20868
rect 4856 20828 4901 20856
rect 5863 20828 5908 20856
rect 4856 20816 4862 20828
rect 5902 20816 5908 20828
rect 5960 20816 5966 20868
rect 5994 20816 6000 20868
rect 6052 20856 6058 20868
rect 6052 20828 6097 20856
rect 6052 20816 6058 20828
rect 7282 20816 7288 20868
rect 7340 20856 7346 20868
rect 7469 20859 7527 20865
rect 7469 20856 7481 20859
rect 7340 20828 7481 20856
rect 7340 20816 7346 20828
rect 7469 20825 7481 20828
rect 7515 20825 7527 20859
rect 7469 20819 7527 20825
rect 7558 20816 7564 20868
rect 7616 20856 7622 20868
rect 8113 20859 8171 20865
rect 7616 20828 7661 20856
rect 7616 20816 7622 20828
rect 8113 20825 8125 20859
rect 8159 20856 8171 20859
rect 8294 20856 8300 20868
rect 8159 20828 8300 20856
rect 8159 20825 8171 20828
rect 8113 20819 8171 20825
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 9214 20816 9220 20868
rect 9272 20856 9278 20868
rect 9324 20856 9352 20887
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 11793 20927 11851 20933
rect 11793 20924 11805 20927
rect 11204 20896 11805 20924
rect 11204 20884 11210 20896
rect 11793 20893 11805 20896
rect 11839 20893 11851 20927
rect 11793 20887 11851 20893
rect 9858 20856 9864 20868
rect 9272 20828 9352 20856
rect 9416 20828 9864 20856
rect 9272 20816 9278 20828
rect 4065 20791 4123 20797
rect 4065 20757 4077 20791
rect 4111 20788 4123 20791
rect 4890 20788 4896 20800
rect 4111 20760 4896 20788
rect 4111 20757 4123 20760
rect 4065 20751 4123 20757
rect 4890 20748 4896 20760
rect 4948 20748 4954 20800
rect 6546 20748 6552 20800
rect 6604 20788 6610 20800
rect 9416 20788 9444 20828
rect 9858 20816 9864 20828
rect 9916 20816 9922 20868
rect 10137 20859 10195 20865
rect 10137 20825 10149 20859
rect 10183 20825 10195 20859
rect 10137 20819 10195 20825
rect 12621 20859 12679 20865
rect 12621 20825 12633 20859
rect 12667 20825 12679 20859
rect 12621 20819 12679 20825
rect 13541 20859 13599 20865
rect 13541 20825 13553 20859
rect 13587 20856 13599 20859
rect 13630 20856 13636 20868
rect 13587 20828 13636 20856
rect 13587 20825 13599 20828
rect 13541 20819 13599 20825
rect 6604 20760 9444 20788
rect 6604 20748 6610 20760
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 10152 20788 10180 20819
rect 9732 20760 10180 20788
rect 11885 20791 11943 20797
rect 9732 20748 9738 20760
rect 11885 20757 11897 20791
rect 11931 20788 11943 20791
rect 12636 20788 12664 20819
rect 13630 20816 13636 20828
rect 13688 20816 13694 20868
rect 14369 20859 14427 20865
rect 14369 20825 14381 20859
rect 14415 20825 14427 20859
rect 14369 20819 14427 20825
rect 14461 20859 14519 20865
rect 14461 20825 14473 20859
rect 14507 20856 14519 20859
rect 14550 20856 14556 20868
rect 14507 20828 14556 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 11931 20760 12664 20788
rect 14384 20788 14412 20819
rect 14550 20816 14556 20828
rect 14608 20816 14614 20868
rect 14734 20816 14740 20868
rect 14792 20856 14798 20868
rect 15120 20856 15148 20964
rect 15194 20884 15200 20936
rect 15252 20924 15258 20936
rect 15657 20927 15715 20933
rect 15657 20924 15669 20927
rect 15252 20896 15669 20924
rect 15252 20884 15258 20896
rect 15657 20893 15669 20896
rect 15703 20893 15715 20927
rect 15764 20924 15792 20964
rect 16942 20952 16948 20964
rect 17000 20952 17006 21004
rect 17218 20992 17224 21004
rect 17131 20964 17224 20992
rect 17218 20952 17224 20964
rect 17276 20992 17282 21004
rect 17402 20992 17408 21004
rect 17276 20964 17408 20992
rect 17276 20952 17282 20964
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 17512 21001 17540 21032
rect 23750 21020 23756 21072
rect 23808 21060 23814 21072
rect 23937 21063 23995 21069
rect 23937 21060 23949 21063
rect 23808 21032 23949 21060
rect 23808 21020 23814 21032
rect 23937 21029 23949 21032
rect 23983 21060 23995 21063
rect 24118 21060 24124 21072
rect 23983 21032 24124 21060
rect 23983 21029 23995 21032
rect 23937 21023 23995 21029
rect 24118 21020 24124 21032
rect 24176 21020 24182 21072
rect 24228 21060 24256 21100
rect 26234 21088 26240 21100
rect 26292 21088 26298 21140
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 29825 21131 29883 21137
rect 29825 21128 29837 21131
rect 26384 21100 29837 21128
rect 26384 21088 26390 21100
rect 29825 21097 29837 21100
rect 29871 21097 29883 21131
rect 29825 21091 29883 21097
rect 32585 21131 32643 21137
rect 32585 21097 32597 21131
rect 32631 21128 32643 21131
rect 36078 21128 36084 21140
rect 32631 21100 36084 21128
rect 32631 21097 32643 21100
rect 32585 21091 32643 21097
rect 36078 21088 36084 21100
rect 36136 21088 36142 21140
rect 24228 21032 26188 21060
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 21784 20964 25544 20992
rect 21784 20952 21790 20964
rect 16206 20924 16212 20936
rect 15764 20896 16212 20924
rect 15657 20887 15715 20893
rect 16206 20884 16212 20896
rect 16264 20884 16270 20936
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 14792 20828 15148 20856
rect 14792 20816 14798 20828
rect 15930 20816 15936 20868
rect 15988 20856 15994 20868
rect 16316 20856 16344 20887
rect 18414 20884 18420 20936
rect 18472 20924 18478 20936
rect 25516 20933 25544 20964
rect 26160 20933 26188 21032
rect 29914 20992 29920 21004
rect 26988 20964 29920 20992
rect 26988 20933 27016 20964
rect 29914 20952 29920 20964
rect 29972 20952 29978 21004
rect 31726 20964 37780 20992
rect 20441 20927 20499 20933
rect 20441 20924 20453 20927
rect 18472 20896 20453 20924
rect 18472 20884 18478 20896
rect 20441 20893 20453 20896
rect 20487 20893 20499 20927
rect 20441 20887 20499 20893
rect 25501 20927 25559 20933
rect 25501 20893 25513 20927
rect 25547 20893 25559 20927
rect 25501 20887 25559 20893
rect 26145 20927 26203 20933
rect 26145 20893 26157 20927
rect 26191 20924 26203 20927
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 26191 20896 26985 20924
rect 26191 20893 26203 20896
rect 26145 20887 26203 20893
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20924 29791 20927
rect 31726 20924 31754 20964
rect 29779 20896 31754 20924
rect 32769 20927 32827 20933
rect 29779 20893 29791 20896
rect 29733 20887 29791 20893
rect 32769 20893 32781 20927
rect 32815 20893 32827 20927
rect 32769 20887 32827 20893
rect 15988 20828 16344 20856
rect 17313 20859 17371 20865
rect 15988 20816 15994 20828
rect 17313 20825 17325 20859
rect 17359 20825 17371 20859
rect 17313 20819 17371 20825
rect 15194 20788 15200 20800
rect 14384 20760 15200 20788
rect 11931 20757 11943 20760
rect 11885 20751 11943 20757
rect 15194 20748 15200 20760
rect 15252 20788 15258 20800
rect 15378 20788 15384 20800
rect 15252 20760 15384 20788
rect 15252 20748 15258 20760
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 15473 20791 15531 20797
rect 15473 20757 15485 20791
rect 15519 20788 15531 20791
rect 15746 20788 15752 20800
rect 15519 20760 15752 20788
rect 15519 20757 15531 20760
rect 15473 20751 15531 20757
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 17328 20788 17356 20819
rect 22370 20816 22376 20868
rect 22428 20856 22434 20868
rect 23385 20859 23443 20865
rect 23385 20856 23397 20859
rect 22428 20828 23397 20856
rect 22428 20816 22434 20828
rect 23385 20825 23397 20828
rect 23431 20825 23443 20859
rect 23385 20819 23443 20825
rect 23477 20859 23535 20865
rect 23477 20825 23489 20859
rect 23523 20856 23535 20859
rect 23842 20856 23848 20868
rect 23523 20828 23848 20856
rect 23523 20825 23535 20828
rect 23477 20819 23535 20825
rect 23842 20816 23848 20828
rect 23900 20816 23906 20868
rect 25593 20859 25651 20865
rect 25593 20825 25605 20859
rect 25639 20856 25651 20859
rect 32784 20856 32812 20887
rect 37182 20884 37188 20936
rect 37240 20924 37246 20936
rect 37752 20933 37780 20964
rect 37461 20927 37519 20933
rect 37461 20924 37473 20927
rect 37240 20896 37473 20924
rect 37240 20884 37246 20896
rect 37461 20893 37473 20896
rect 37507 20893 37519 20927
rect 37461 20887 37519 20893
rect 37737 20927 37795 20933
rect 37737 20893 37749 20927
rect 37783 20924 37795 20927
rect 37826 20924 37832 20936
rect 37783 20896 37832 20924
rect 37783 20893 37795 20896
rect 37737 20887 37795 20893
rect 37826 20884 37832 20896
rect 37884 20884 37890 20936
rect 25639 20828 32812 20856
rect 25639 20825 25651 20828
rect 25593 20819 25651 20825
rect 18138 20788 18144 20800
rect 17328 20760 18144 20788
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 24854 20788 24860 20800
rect 24815 20760 24860 20788
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 26786 20788 26792 20800
rect 26747 20760 26792 20788
rect 26786 20748 26792 20760
rect 26844 20748 26850 20800
rect 29914 20748 29920 20800
rect 29972 20788 29978 20800
rect 37734 20788 37740 20800
rect 29972 20760 37740 20788
rect 29972 20748 29978 20760
rect 37734 20748 37740 20760
rect 37792 20748 37798 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1302 20544 1308 20596
rect 1360 20584 1366 20596
rect 2038 20584 2044 20596
rect 1360 20556 2044 20584
rect 1360 20544 1366 20556
rect 2038 20544 2044 20556
rect 2096 20544 2102 20596
rect 4430 20584 4436 20596
rect 3344 20556 4436 20584
rect 1670 20516 1676 20528
rect 1631 20488 1676 20516
rect 1670 20476 1676 20488
rect 1728 20476 1734 20528
rect 1765 20519 1823 20525
rect 1765 20485 1777 20519
rect 1811 20516 1823 20519
rect 1946 20516 1952 20528
rect 1811 20488 1952 20516
rect 1811 20485 1823 20488
rect 1765 20479 1823 20485
rect 1946 20476 1952 20488
rect 2004 20476 2010 20528
rect 2590 20476 2596 20528
rect 2648 20516 2654 20528
rect 3344 20525 3372 20556
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4982 20544 4988 20596
rect 5040 20544 5046 20596
rect 7926 20584 7932 20596
rect 5092 20556 7932 20584
rect 2685 20519 2743 20525
rect 2685 20516 2697 20519
rect 2648 20488 2697 20516
rect 2648 20476 2654 20488
rect 2685 20485 2697 20488
rect 2731 20485 2743 20519
rect 2685 20479 2743 20485
rect 3329 20519 3387 20525
rect 3329 20485 3341 20519
rect 3375 20485 3387 20519
rect 3329 20479 3387 20485
rect 3881 20519 3939 20525
rect 3881 20485 3893 20519
rect 3927 20516 3939 20519
rect 3970 20516 3976 20528
rect 3927 20488 3976 20516
rect 3927 20485 3939 20488
rect 3881 20479 3939 20485
rect 3970 20476 3976 20488
rect 4028 20476 4034 20528
rect 4525 20519 4583 20525
rect 4525 20485 4537 20519
rect 4571 20516 4583 20519
rect 5000 20516 5028 20544
rect 5092 20525 5120 20556
rect 7926 20544 7932 20556
rect 7984 20544 7990 20596
rect 8846 20544 8852 20596
rect 8904 20584 8910 20596
rect 11238 20584 11244 20596
rect 8904 20556 10364 20584
rect 8904 20544 8910 20556
rect 4571 20488 5028 20516
rect 5077 20519 5135 20525
rect 4571 20485 4583 20488
rect 4525 20479 4583 20485
rect 5077 20485 5089 20519
rect 5123 20485 5135 20519
rect 6638 20516 6644 20528
rect 6599 20488 6644 20516
rect 5077 20479 5135 20485
rect 6638 20476 6644 20488
rect 6696 20476 6702 20528
rect 6733 20519 6791 20525
rect 6733 20485 6745 20519
rect 6779 20516 6791 20519
rect 7098 20516 7104 20528
rect 6779 20488 7104 20516
rect 6779 20485 6791 20488
rect 6733 20479 6791 20485
rect 7098 20476 7104 20488
rect 7156 20476 7162 20528
rect 8205 20519 8263 20525
rect 8205 20485 8217 20519
rect 8251 20516 8263 20519
rect 8754 20516 8760 20528
rect 8251 20488 8760 20516
rect 8251 20485 8263 20488
rect 8205 20479 8263 20485
rect 8754 20476 8760 20488
rect 8812 20476 8818 20528
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 5994 20448 6000 20460
rect 5859 20420 6000 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 3237 20383 3295 20389
rect 3237 20349 3249 20383
rect 3283 20380 3295 20383
rect 3326 20380 3332 20392
rect 3283 20352 3332 20380
rect 3283 20349 3295 20352
rect 3237 20343 3295 20349
rect 3326 20340 3332 20352
rect 3384 20340 3390 20392
rect 4433 20383 4491 20389
rect 4433 20349 4445 20383
rect 4479 20380 4491 20383
rect 5902 20380 5908 20392
rect 4479 20352 5908 20380
rect 4479 20349 4491 20352
rect 4433 20343 4491 20349
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 6914 20380 6920 20392
rect 6875 20352 6920 20380
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 9030 20380 9036 20392
rect 8159 20352 9036 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 9125 20383 9183 20389
rect 9125 20349 9137 20383
rect 9171 20349 9183 20383
rect 9766 20380 9772 20392
rect 9727 20352 9772 20380
rect 9125 20343 9183 20349
rect 4706 20272 4712 20324
rect 4764 20312 4770 20324
rect 6178 20312 6184 20324
rect 4764 20284 6184 20312
rect 4764 20272 4770 20284
rect 6178 20272 6184 20284
rect 6236 20272 6242 20324
rect 6638 20272 6644 20324
rect 6696 20312 6702 20324
rect 9140 20312 9168 20343
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 10336 20380 10364 20556
rect 10612 20556 11244 20584
rect 10502 20516 10508 20528
rect 10463 20488 10508 20516
rect 10502 20476 10508 20488
rect 10560 20476 10566 20528
rect 10612 20525 10640 20556
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 12584 20556 12664 20584
rect 12584 20544 12590 20556
rect 10597 20519 10655 20525
rect 10597 20485 10609 20519
rect 10643 20485 10655 20519
rect 10597 20479 10655 20485
rect 10870 20476 10876 20528
rect 10928 20516 10934 20528
rect 11885 20519 11943 20525
rect 11885 20516 11897 20519
rect 10928 20488 11897 20516
rect 10928 20476 10934 20488
rect 11885 20485 11897 20488
rect 11931 20485 11943 20519
rect 11885 20479 11943 20485
rect 12636 20392 12664 20556
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 17589 20587 17647 20593
rect 13688 20556 16528 20584
rect 13688 20544 13694 20556
rect 12805 20519 12863 20525
rect 12805 20485 12817 20519
rect 12851 20516 12863 20519
rect 13170 20516 13176 20528
rect 12851 20488 13176 20516
rect 12851 20485 12863 20488
rect 12805 20479 12863 20485
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 14844 20525 14872 20556
rect 13806 20519 13864 20525
rect 13806 20516 13818 20519
rect 13596 20488 13818 20516
rect 13596 20476 13602 20488
rect 13806 20485 13818 20488
rect 13852 20485 13864 20519
rect 13806 20479 13864 20485
rect 13918 20519 13976 20525
rect 13918 20485 13930 20519
rect 13964 20516 13976 20519
rect 14829 20519 14887 20525
rect 13964 20488 14780 20516
rect 13964 20485 13976 20488
rect 13918 20479 13976 20485
rect 14752 20448 14780 20488
rect 14829 20485 14841 20519
rect 14875 20485 14887 20519
rect 15470 20516 15476 20528
rect 15431 20488 15476 20516
rect 14829 20479 14887 20485
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 15102 20448 15108 20460
rect 14752 20420 15108 20448
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 11793 20383 11851 20389
rect 11793 20380 11805 20383
rect 10336 20368 10732 20380
rect 10888 20368 11805 20380
rect 10336 20352 11805 20368
rect 10704 20340 10916 20352
rect 11793 20349 11805 20352
rect 11839 20349 11851 20383
rect 11793 20343 11851 20349
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 15381 20383 15439 20389
rect 15381 20349 15393 20383
rect 15427 20349 15439 20383
rect 15654 20380 15660 20392
rect 15615 20352 15660 20380
rect 15381 20343 15439 20349
rect 6696 20284 6868 20312
rect 9140 20284 9352 20312
rect 6696 20272 6702 20284
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 6730 20244 6736 20256
rect 5951 20216 6736 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 6840 20244 6868 20284
rect 7006 20244 7012 20256
rect 6840 20216 7012 20244
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9122 20244 9128 20256
rect 8352 20216 9128 20244
rect 8352 20204 8358 20216
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 9324 20244 9352 20284
rect 9490 20272 9496 20324
rect 9548 20312 9554 20324
rect 11057 20315 11115 20321
rect 11057 20312 11069 20315
rect 9548 20284 11069 20312
rect 9548 20272 9554 20284
rect 11057 20281 11069 20284
rect 11103 20281 11115 20315
rect 11057 20275 11115 20281
rect 10870 20244 10876 20256
rect 9324 20216 10876 20244
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 11072 20244 11100 20275
rect 12894 20272 12900 20324
rect 12952 20312 12958 20324
rect 13446 20312 13452 20324
rect 12952 20284 13452 20312
rect 12952 20272 12958 20284
rect 13446 20272 13452 20284
rect 13504 20312 13510 20324
rect 15396 20312 15424 20343
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 13504 20284 15424 20312
rect 16500 20312 16528 20556
rect 17589 20553 17601 20587
rect 17635 20584 17647 20587
rect 22370 20584 22376 20596
rect 17635 20556 22376 20584
rect 17635 20553 17647 20556
rect 17589 20547 17647 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 23658 20584 23664 20596
rect 23619 20556 23664 20584
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 23842 20544 23848 20596
rect 23900 20584 23906 20596
rect 24213 20587 24271 20593
rect 24213 20584 24225 20587
rect 23900 20556 24225 20584
rect 23900 20544 23906 20556
rect 24213 20553 24225 20556
rect 24259 20553 24271 20587
rect 26694 20584 26700 20596
rect 24213 20547 24271 20553
rect 24320 20556 26700 20584
rect 17218 20476 17224 20528
rect 17276 20516 17282 20528
rect 18509 20519 18567 20525
rect 18509 20516 18521 20519
rect 17276 20488 18521 20516
rect 17276 20476 17282 20488
rect 18509 20485 18521 20488
rect 18555 20485 18567 20519
rect 24320 20516 24348 20556
rect 26694 20544 26700 20556
rect 26752 20544 26758 20596
rect 25774 20516 25780 20528
rect 18509 20479 18567 20485
rect 22066 20488 24348 20516
rect 25735 20488 25780 20516
rect 16942 20448 16948 20460
rect 16903 20420 16948 20448
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20448 17187 20451
rect 17954 20448 17960 20460
rect 17175 20420 17960 20448
rect 17175 20417 17187 20420
rect 17129 20411 17187 20417
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 22066 20448 22094 20488
rect 25774 20476 25780 20488
rect 25832 20476 25838 20528
rect 23566 20448 23572 20460
rect 19352 20420 22094 20448
rect 23527 20420 23572 20448
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 18417 20383 18475 20389
rect 18417 20380 18429 20383
rect 17920 20352 18429 20380
rect 17920 20340 17926 20352
rect 18417 20349 18429 20352
rect 18463 20380 18475 20383
rect 19352 20380 19380 20420
rect 23566 20408 23572 20420
rect 23624 20408 23630 20460
rect 24394 20448 24400 20460
rect 24355 20420 24400 20448
rect 24394 20408 24400 20420
rect 24452 20408 24458 20460
rect 18463 20352 19380 20380
rect 19429 20383 19487 20389
rect 18463 20349 18475 20352
rect 18417 20343 18475 20349
rect 19429 20349 19441 20383
rect 19475 20349 19487 20383
rect 19429 20343 19487 20349
rect 19058 20312 19064 20324
rect 16500 20284 19064 20312
rect 13504 20272 13510 20284
rect 19058 20272 19064 20284
rect 19116 20312 19122 20324
rect 19444 20312 19472 20343
rect 24854 20340 24860 20392
rect 24912 20380 24918 20392
rect 25685 20383 25743 20389
rect 25685 20380 25697 20383
rect 24912 20352 25697 20380
rect 24912 20340 24918 20352
rect 25685 20349 25697 20352
rect 25731 20349 25743 20383
rect 25685 20343 25743 20349
rect 26329 20383 26387 20389
rect 26329 20349 26341 20383
rect 26375 20380 26387 20383
rect 26510 20380 26516 20392
rect 26375 20352 26516 20380
rect 26375 20349 26387 20352
rect 26329 20343 26387 20349
rect 26510 20340 26516 20352
rect 26568 20380 26574 20392
rect 26970 20380 26976 20392
rect 26568 20352 26976 20380
rect 26568 20340 26574 20352
rect 26970 20340 26976 20352
rect 27028 20340 27034 20392
rect 19116 20284 19472 20312
rect 19116 20272 19122 20284
rect 19518 20272 19524 20324
rect 19576 20312 19582 20324
rect 22554 20312 22560 20324
rect 19576 20284 22560 20312
rect 19576 20272 19582 20284
rect 22554 20272 22560 20284
rect 22612 20272 22618 20324
rect 17310 20244 17316 20256
rect 11072 20216 17316 20244
rect 17310 20204 17316 20216
rect 17368 20204 17374 20256
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 26878 20244 26884 20256
rect 18932 20216 26884 20244
rect 18932 20204 18938 20216
rect 26878 20204 26884 20216
rect 26936 20204 26942 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 4798 20000 4804 20052
rect 4856 20040 4862 20052
rect 4856 20012 9628 20040
rect 4856 20000 4862 20012
rect 6914 19972 6920 19984
rect 2424 19944 6920 19972
rect 2424 19913 2452 19944
rect 6914 19932 6920 19944
rect 6972 19972 6978 19984
rect 9490 19972 9496 19984
rect 6972 19944 9496 19972
rect 6972 19932 6978 19944
rect 9490 19932 9496 19944
rect 9548 19932 9554 19984
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 4706 19904 4712 19916
rect 3467 19876 4712 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 4706 19864 4712 19876
rect 4764 19864 4770 19916
rect 4798 19864 4804 19916
rect 4856 19904 4862 19916
rect 5077 19907 5135 19913
rect 5077 19904 5089 19907
rect 4856 19876 5089 19904
rect 4856 19864 4862 19876
rect 5077 19873 5089 19876
rect 5123 19873 5135 19907
rect 5077 19867 5135 19873
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 7837 19907 7895 19913
rect 7837 19904 7849 19907
rect 6236 19876 7849 19904
rect 6236 19864 6242 19876
rect 7837 19873 7849 19876
rect 7883 19904 7895 19907
rect 8386 19904 8392 19916
rect 7883 19876 8392 19904
rect 7883 19873 7895 19876
rect 7837 19867 7895 19873
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 9600 19913 9628 20012
rect 10870 20000 10876 20052
rect 10928 20040 10934 20052
rect 15378 20040 15384 20052
rect 10928 20012 15384 20040
rect 10928 20000 10934 20012
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 16390 20040 16396 20052
rect 16351 20012 16396 20040
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 18138 20040 18144 20052
rect 18099 20012 18144 20040
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 25774 20040 25780 20052
rect 18380 20012 22600 20040
rect 25735 20012 25780 20040
rect 18380 20000 18386 20012
rect 13170 19932 13176 19984
rect 13228 19972 13234 19984
rect 13814 19972 13820 19984
rect 13228 19944 13820 19972
rect 13228 19932 13234 19944
rect 13814 19932 13820 19944
rect 13872 19932 13878 19984
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 21634 19972 21640 19984
rect 17184 19944 21640 19972
rect 17184 19932 17190 19944
rect 21634 19932 21640 19944
rect 21692 19932 21698 19984
rect 9585 19907 9643 19913
rect 9585 19873 9597 19907
rect 9631 19873 9643 19907
rect 9585 19867 9643 19873
rect 9766 19864 9772 19916
rect 9824 19904 9830 19916
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 9824 19876 10517 19904
rect 9824 19864 9830 19876
rect 10505 19873 10517 19876
rect 10551 19873 10563 19907
rect 12066 19904 12072 19916
rect 12027 19876 12072 19904
rect 10505 19867 10563 19873
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 13538 19904 13544 19916
rect 13499 19876 13544 19904
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 14369 19907 14427 19913
rect 14369 19873 14381 19907
rect 14415 19904 14427 19907
rect 16666 19904 16672 19916
rect 14415 19876 16672 19904
rect 14415 19873 14427 19876
rect 14369 19867 14427 19873
rect 16666 19864 16672 19876
rect 16724 19864 16730 19916
rect 17310 19864 17316 19916
rect 17368 19904 17374 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 17368 19876 21741 19904
rect 17368 19864 17374 19876
rect 21729 19873 21741 19876
rect 21775 19873 21787 19907
rect 21729 19867 21787 19873
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 1854 19836 1860 19848
rect 1811 19808 1860 19836
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 4338 19836 4344 19848
rect 4299 19808 4344 19836
rect 4338 19796 4344 19808
rect 4396 19796 4402 19848
rect 6546 19796 6552 19848
rect 6604 19836 6610 19848
rect 6825 19839 6883 19845
rect 6825 19836 6837 19839
rect 6604 19808 6837 19836
rect 6604 19796 6610 19808
rect 6825 19805 6837 19808
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 15746 19796 15752 19848
rect 15804 19836 15810 19848
rect 16301 19839 16359 19845
rect 16301 19836 16313 19839
rect 15804 19808 16313 19836
rect 15804 19796 15810 19808
rect 16301 19805 16313 19808
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19838 17095 19839
rect 17083 19836 17172 19838
rect 17494 19836 17500 19848
rect 17083 19810 17500 19836
rect 17083 19805 17095 19810
rect 17144 19808 17500 19810
rect 17037 19799 17095 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19838 18107 19839
rect 18095 19810 18184 19838
rect 18095 19805 18107 19810
rect 18049 19799 18107 19805
rect 18156 19780 18184 19810
rect 18598 19796 18604 19848
rect 18656 19836 18662 19848
rect 19518 19836 19524 19848
rect 18656 19808 19524 19836
rect 18656 19796 18662 19808
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 22572 19845 22600 20012
rect 25774 20000 25780 20012
rect 25832 20000 25838 20052
rect 25498 19972 25504 19984
rect 23216 19944 25504 19972
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 2498 19728 2504 19780
rect 2556 19768 2562 19780
rect 2556 19740 2601 19768
rect 2556 19728 2562 19740
rect 5166 19728 5172 19780
rect 5224 19768 5230 19780
rect 6089 19771 6147 19777
rect 5224 19740 5269 19768
rect 5224 19728 5230 19740
rect 6089 19737 6101 19771
rect 6135 19768 6147 19771
rect 6178 19768 6184 19780
rect 6135 19740 6184 19768
rect 6135 19737 6147 19740
rect 6089 19731 6147 19737
rect 6178 19728 6184 19740
rect 6236 19728 6242 19780
rect 7006 19768 7012 19780
rect 6967 19740 7012 19768
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 7561 19771 7619 19777
rect 7561 19737 7573 19771
rect 7607 19737 7619 19771
rect 7561 19731 7619 19737
rect 1765 19703 1823 19709
rect 1765 19669 1777 19703
rect 1811 19700 1823 19703
rect 3694 19700 3700 19712
rect 1811 19672 3700 19700
rect 1811 19669 1823 19672
rect 1765 19663 1823 19669
rect 3694 19660 3700 19672
rect 3752 19660 3758 19712
rect 4433 19703 4491 19709
rect 4433 19669 4445 19703
rect 4479 19700 4491 19703
rect 4706 19700 4712 19712
rect 4479 19672 4712 19700
rect 4479 19669 4491 19672
rect 4433 19663 4491 19669
rect 4706 19660 4712 19672
rect 4764 19660 4770 19712
rect 7576 19700 7604 19731
rect 7650 19728 7656 19780
rect 7708 19768 7714 19780
rect 9309 19771 9367 19777
rect 7708 19740 7753 19768
rect 7708 19728 7714 19740
rect 9309 19737 9321 19771
rect 9355 19737 9367 19771
rect 9309 19731 9367 19737
rect 8938 19700 8944 19712
rect 7576 19672 8944 19700
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 9324 19700 9352 19731
rect 9398 19728 9404 19780
rect 9456 19768 9462 19780
rect 9456 19740 9501 19768
rect 9456 19728 9462 19740
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 10597 19771 10655 19777
rect 10597 19768 10609 19771
rect 10192 19740 10609 19768
rect 10192 19728 10198 19740
rect 10597 19737 10609 19740
rect 10643 19737 10655 19771
rect 11514 19768 11520 19780
rect 11475 19740 11520 19768
rect 10597 19731 10655 19737
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 12158 19768 12164 19780
rect 12119 19740 12164 19768
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 13081 19771 13139 19777
rect 13081 19737 13093 19771
rect 13127 19768 13139 19771
rect 13170 19768 13176 19780
rect 13127 19740 13176 19768
rect 13127 19737 13139 19740
rect 13081 19731 13139 19737
rect 13170 19728 13176 19740
rect 13228 19728 13234 19780
rect 14458 19728 14464 19780
rect 14516 19768 14522 19780
rect 15378 19768 15384 19780
rect 14516 19740 14561 19768
rect 15339 19740 15384 19768
rect 14516 19728 14522 19740
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 16592 19740 18000 19768
rect 12710 19700 12716 19712
rect 9324 19672 12716 19700
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 16592 19700 16620 19740
rect 14240 19672 16620 19700
rect 14240 19660 14246 19672
rect 16666 19660 16672 19712
rect 16724 19700 16730 19712
rect 17129 19703 17187 19709
rect 17129 19700 17141 19703
rect 16724 19672 17141 19700
rect 16724 19660 16730 19672
rect 17129 19669 17141 19672
rect 17175 19669 17187 19703
rect 17972 19700 18000 19740
rect 18138 19728 18144 19780
rect 18196 19728 18202 19780
rect 20346 19768 20352 19780
rect 18248 19740 20352 19768
rect 18248 19700 18276 19740
rect 20346 19728 20352 19740
rect 20404 19728 20410 19780
rect 21450 19768 21456 19780
rect 21411 19740 21456 19768
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 21545 19771 21603 19777
rect 21545 19737 21557 19771
rect 21591 19737 21603 19771
rect 21545 19731 21603 19737
rect 17972 19672 18276 19700
rect 21560 19700 21588 19731
rect 21634 19728 21640 19780
rect 21692 19768 21698 19780
rect 23216 19768 23244 19944
rect 25498 19932 25504 19944
rect 25556 19932 25562 19984
rect 23382 19904 23388 19916
rect 23343 19876 23388 19904
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 24026 19904 24032 19916
rect 23987 19876 24032 19904
rect 24026 19864 24032 19876
rect 24084 19864 24090 19916
rect 26878 19864 26884 19916
rect 26936 19904 26942 19916
rect 35526 19904 35532 19916
rect 26936 19876 35532 19904
rect 26936 19864 26942 19876
rect 35526 19864 35532 19876
rect 35584 19864 35590 19916
rect 24578 19836 24584 19848
rect 24539 19808 24584 19836
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19836 26019 19839
rect 26786 19836 26792 19848
rect 26007 19808 26792 19836
rect 26007 19805 26019 19808
rect 25961 19799 26019 19805
rect 26786 19796 26792 19808
rect 26844 19796 26850 19848
rect 26970 19796 26976 19848
rect 27028 19836 27034 19848
rect 32033 19839 32091 19845
rect 32033 19836 32045 19839
rect 27028 19808 32045 19836
rect 27028 19796 27034 19808
rect 32033 19805 32045 19808
rect 32079 19805 32091 19839
rect 32033 19799 32091 19805
rect 21692 19740 23244 19768
rect 23477 19771 23535 19777
rect 21692 19728 21698 19740
rect 23477 19737 23489 19771
rect 23523 19768 23535 19771
rect 23523 19740 23704 19768
rect 23523 19737 23535 19740
rect 23477 19731 23535 19737
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 21560 19672 22661 19700
rect 17129 19663 17187 19669
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 23676 19700 23704 19740
rect 23934 19700 23940 19712
rect 23676 19672 23940 19700
rect 22649 19663 22707 19669
rect 23934 19660 23940 19672
rect 23992 19660 23998 19712
rect 24673 19703 24731 19709
rect 24673 19669 24685 19703
rect 24719 19700 24731 19703
rect 24946 19700 24952 19712
rect 24719 19672 24952 19700
rect 24719 19669 24731 19672
rect 24673 19663 24731 19669
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 32125 19703 32183 19709
rect 32125 19669 32137 19703
rect 32171 19700 32183 19703
rect 34422 19700 34428 19712
rect 32171 19672 34428 19700
rect 32171 19669 32183 19672
rect 32125 19663 32183 19669
rect 34422 19660 34428 19672
rect 34480 19660 34486 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3694 19496 3700 19508
rect 1688 19468 3700 19496
rect 1688 19437 1716 19468
rect 3694 19456 3700 19468
rect 3752 19496 3758 19508
rect 6825 19499 6883 19505
rect 3752 19468 6776 19496
rect 3752 19456 3758 19468
rect 1673 19431 1731 19437
rect 1673 19397 1685 19431
rect 1719 19397 1731 19431
rect 1673 19391 1731 19397
rect 1765 19431 1823 19437
rect 1765 19397 1777 19431
rect 1811 19428 1823 19431
rect 2130 19428 2136 19440
rect 1811 19400 2136 19428
rect 1811 19397 1823 19400
rect 1765 19391 1823 19397
rect 2130 19388 2136 19400
rect 2188 19388 2194 19440
rect 2590 19388 2596 19440
rect 2648 19428 2654 19440
rect 2685 19431 2743 19437
rect 2685 19428 2697 19431
rect 2648 19400 2697 19428
rect 2648 19388 2654 19400
rect 2685 19397 2697 19400
rect 2731 19397 2743 19431
rect 2685 19391 2743 19397
rect 5258 19388 5264 19440
rect 5316 19388 5322 19440
rect 6748 19428 6776 19468
rect 6825 19465 6837 19499
rect 6871 19496 6883 19499
rect 6871 19468 10272 19496
rect 6871 19465 6883 19468
rect 6825 19459 6883 19465
rect 7282 19428 7288 19440
rect 6748 19400 7288 19428
rect 7282 19388 7288 19400
rect 7340 19388 7346 19440
rect 9950 19428 9956 19440
rect 8878 19400 9956 19428
rect 9950 19388 9956 19400
rect 10008 19388 10014 19440
rect 10244 19437 10272 19468
rect 10962 19456 10968 19508
rect 11020 19496 11026 19508
rect 14918 19496 14924 19508
rect 11020 19468 14924 19496
rect 11020 19456 11026 19468
rect 14918 19456 14924 19468
rect 14976 19456 14982 19508
rect 15102 19456 15108 19508
rect 15160 19496 15166 19508
rect 16945 19499 17003 19505
rect 16945 19496 16957 19499
rect 15160 19468 16957 19496
rect 15160 19456 15166 19468
rect 16945 19465 16957 19468
rect 16991 19465 17003 19499
rect 16945 19459 17003 19465
rect 21450 19456 21456 19508
rect 21508 19496 21514 19508
rect 23934 19496 23940 19508
rect 21508 19468 23520 19496
rect 23895 19468 23940 19496
rect 21508 19456 21514 19468
rect 10229 19431 10287 19437
rect 10229 19397 10241 19431
rect 10275 19397 10287 19431
rect 10229 19391 10287 19397
rect 12161 19431 12219 19437
rect 12161 19397 12173 19431
rect 12207 19428 12219 19431
rect 12897 19431 12955 19437
rect 12897 19428 12909 19431
rect 12207 19400 12909 19428
rect 12207 19397 12219 19400
rect 12161 19391 12219 19397
rect 12897 19397 12909 19400
rect 12943 19397 12955 19431
rect 14182 19428 14188 19440
rect 14143 19400 14188 19428
rect 12897 19391 12955 19397
rect 14182 19388 14188 19400
rect 14240 19388 14246 19440
rect 14277 19431 14335 19437
rect 14277 19397 14289 19431
rect 14323 19428 14335 19431
rect 15749 19431 15807 19437
rect 15749 19428 15761 19431
rect 14323 19400 15761 19428
rect 14323 19397 14335 19400
rect 14277 19391 14335 19397
rect 15749 19397 15761 19400
rect 15795 19397 15807 19431
rect 15749 19391 15807 19397
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 17957 19431 18015 19437
rect 17957 19428 17969 19431
rect 16632 19400 17969 19428
rect 16632 19388 16638 19400
rect 17957 19397 17969 19400
rect 18003 19397 18015 19431
rect 17957 19391 18015 19397
rect 18138 19388 18144 19440
rect 18196 19428 18202 19440
rect 18322 19428 18328 19440
rect 18196 19400 18328 19428
rect 18196 19388 18202 19400
rect 18322 19388 18328 19400
rect 18380 19388 18386 19440
rect 18874 19428 18880 19440
rect 18835 19400 18880 19428
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 20073 19431 20131 19437
rect 20073 19397 20085 19431
rect 20119 19428 20131 19431
rect 20254 19428 20260 19440
rect 20119 19400 20260 19428
rect 20119 19397 20131 19400
rect 20073 19391 20131 19397
rect 20254 19388 20260 19400
rect 20312 19428 20318 19440
rect 20622 19428 20628 19440
rect 20312 19400 20628 19428
rect 20312 19388 20318 19400
rect 20622 19388 20628 19400
rect 20680 19388 20686 19440
rect 23492 19428 23520 19468
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 30009 19499 30067 19505
rect 30009 19496 30021 19499
rect 24780 19468 30021 19496
rect 24780 19428 24808 19468
rect 30009 19465 30021 19468
rect 30055 19465 30067 19499
rect 38105 19499 38163 19505
rect 38105 19496 38117 19499
rect 30009 19459 30067 19465
rect 35866 19468 38117 19496
rect 24946 19428 24952 19440
rect 20732 19400 23428 19428
rect 23492 19400 24808 19428
rect 24907 19400 24952 19428
rect 3234 19360 3240 19372
rect 3195 19332 3240 19360
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3970 19360 3976 19372
rect 3931 19332 3976 19360
rect 3970 19320 3976 19332
rect 4028 19320 4034 19372
rect 6733 19363 6791 19369
rect 6733 19360 6745 19363
rect 5552 19332 6745 19360
rect 4706 19252 4712 19304
rect 4764 19292 4770 19304
rect 4982 19292 4988 19304
rect 4764 19264 4988 19292
rect 4764 19252 4770 19264
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 5258 19184 5264 19236
rect 5316 19224 5322 19236
rect 5552 19224 5580 19332
rect 6733 19329 6745 19332
rect 6779 19329 6791 19363
rect 11422 19360 11428 19372
rect 6733 19323 6791 19329
rect 10980 19332 11428 19360
rect 5718 19292 5724 19304
rect 5679 19264 5724 19292
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 6972 19264 7389 19292
rect 6972 19252 6978 19264
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7377 19255 7435 19261
rect 7653 19295 7711 19301
rect 7653 19261 7665 19295
rect 7699 19292 7711 19295
rect 10137 19295 10195 19301
rect 7699 19264 9674 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 9646 19224 9674 19264
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 10226 19292 10232 19304
rect 10183 19264 10232 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10226 19252 10232 19264
rect 10284 19292 10290 19304
rect 10980 19292 11008 19332
rect 11422 19320 11428 19332
rect 11480 19320 11486 19372
rect 12069 19363 12127 19369
rect 12069 19329 12081 19363
rect 12115 19360 12127 19363
rect 12618 19360 12624 19372
rect 12115 19332 12624 19360
rect 12115 19329 12127 19332
rect 12069 19323 12127 19329
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 15102 19320 15108 19372
rect 15160 19360 15166 19372
rect 15654 19360 15660 19372
rect 15160 19332 15516 19360
rect 15615 19332 15660 19360
rect 15160 19320 15166 19332
rect 10284 19264 11008 19292
rect 10284 19252 10290 19264
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 12805 19295 12863 19301
rect 11112 19264 12756 19292
rect 11112 19252 11118 19264
rect 10962 19224 10968 19236
rect 5316 19196 5580 19224
rect 5644 19196 6408 19224
rect 9646 19196 10968 19224
rect 5316 19184 5322 19196
rect 3326 19156 3332 19168
rect 3287 19128 3332 19156
rect 3326 19116 3332 19128
rect 3384 19116 3390 19168
rect 4236 19159 4294 19165
rect 4236 19125 4248 19159
rect 4282 19156 4294 19159
rect 5644 19156 5672 19196
rect 4282 19128 5672 19156
rect 6380 19156 6408 19196
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 12728 19224 12756 19264
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 12894 19292 12900 19304
rect 12851 19264 12900 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 12986 19252 12992 19304
rect 13044 19292 13050 19304
rect 13449 19295 13507 19301
rect 13449 19292 13461 19295
rect 13044 19264 13461 19292
rect 13044 19252 13050 19264
rect 13449 19261 13461 19264
rect 13495 19292 13507 19295
rect 13538 19292 13544 19304
rect 13495 19264 13544 19292
rect 13495 19261 13507 19264
rect 13449 19255 13507 19261
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 14645 19295 14703 19301
rect 14645 19261 14657 19295
rect 14691 19261 14703 19295
rect 15488 19292 15516 19332
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 15764 19332 16865 19360
rect 15764 19292 15792 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 20732 19360 20760 19400
rect 19392 19332 20760 19360
rect 21453 19363 21511 19369
rect 19392 19320 19398 19332
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 22186 19360 22192 19372
rect 21499 19332 22048 19360
rect 22147 19332 22192 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 17862 19292 17868 19304
rect 15488 19264 15792 19292
rect 17823 19264 17868 19292
rect 14645 19255 14703 19261
rect 13170 19224 13176 19236
rect 12728 19196 13176 19224
rect 13170 19184 13176 19196
rect 13228 19224 13234 19236
rect 14660 19224 14688 19255
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 13228 19196 14688 19224
rect 13228 19184 13234 19196
rect 15286 19184 15292 19236
rect 15344 19224 15350 19236
rect 15838 19224 15844 19236
rect 15344 19196 15844 19224
rect 15344 19184 15350 19196
rect 15838 19184 15844 19196
rect 15896 19224 15902 19236
rect 21910 19224 21916 19236
rect 15896 19196 21916 19224
rect 15896 19184 15902 19196
rect 21910 19184 21916 19196
rect 21968 19184 21974 19236
rect 22020 19233 22048 19332
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 23400 19369 23428 19400
rect 24946 19388 24952 19400
rect 25004 19388 25010 19440
rect 25498 19428 25504 19440
rect 25459 19400 25504 19428
rect 25498 19388 25504 19400
rect 25556 19388 25562 19440
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19360 23443 19363
rect 23845 19363 23903 19369
rect 23845 19360 23857 19363
rect 23431 19332 23857 19360
rect 23431 19329 23443 19332
rect 23385 19323 23443 19329
rect 23845 19329 23857 19332
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 29917 19363 29975 19369
rect 29917 19329 29929 19363
rect 29963 19360 29975 19363
rect 35866 19360 35894 19468
rect 38105 19465 38117 19468
rect 38151 19465 38163 19499
rect 38105 19459 38163 19465
rect 38286 19360 38292 19372
rect 29963 19332 35894 19360
rect 38247 19332 38292 19360
rect 29963 19329 29975 19332
rect 29917 19323 29975 19329
rect 38286 19320 38292 19332
rect 38344 19320 38350 19372
rect 24854 19292 24860 19304
rect 24815 19264 24860 19292
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 24946 19252 24952 19304
rect 25004 19292 25010 19304
rect 25961 19295 26019 19301
rect 25961 19292 25973 19295
rect 25004 19264 25973 19292
rect 25004 19252 25010 19264
rect 25961 19261 25973 19264
rect 26007 19261 26019 19295
rect 25961 19255 26019 19261
rect 22005 19227 22063 19233
rect 22005 19193 22017 19227
rect 22051 19193 22063 19227
rect 22005 19187 22063 19193
rect 8018 19156 8024 19168
rect 6380 19128 8024 19156
rect 4282 19125 4294 19128
rect 4236 19119 4294 19125
rect 8018 19116 8024 19128
rect 8076 19116 8082 19168
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 9125 19159 9183 19165
rect 9125 19156 9137 19159
rect 8444 19128 9137 19156
rect 8444 19116 8450 19128
rect 9125 19125 9137 19128
rect 9171 19125 9183 19159
rect 9125 19119 9183 19125
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 12526 19156 12532 19168
rect 9364 19128 12532 19156
rect 9364 19116 9370 19128
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 13780 19128 20177 19156
rect 13780 19116 13786 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 20165 19119 20223 19125
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 23201 19159 23259 19165
rect 23201 19125 23213 19159
rect 23247 19156 23259 19159
rect 23382 19156 23388 19168
rect 23247 19128 23388 19156
rect 23247 19125 23259 19128
rect 23201 19119 23259 19125
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 3329 18955 3387 18961
rect 3329 18921 3341 18955
rect 3375 18952 3387 18955
rect 3418 18952 3424 18964
rect 3375 18924 3424 18952
rect 3375 18921 3387 18924
rect 3329 18915 3387 18921
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 3973 18955 4031 18961
rect 3973 18921 3985 18955
rect 4019 18952 4031 18955
rect 8570 18952 8576 18964
rect 4019 18924 8156 18952
rect 8531 18924 8576 18952
rect 4019 18921 4031 18924
rect 3973 18915 4031 18921
rect 3988 18884 4016 18915
rect 3252 18856 4016 18884
rect 8128 18884 8156 18924
rect 8570 18912 8576 18924
rect 8628 18912 8634 18964
rect 8662 18912 8668 18964
rect 8720 18952 8726 18964
rect 9950 18952 9956 18964
rect 8720 18924 9956 18952
rect 8720 18912 8726 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 15562 18952 15568 18964
rect 15523 18924 15568 18952
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 17218 18952 17224 18964
rect 17179 18924 17224 18952
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19484 18924 19717 18952
rect 19484 18912 19490 18924
rect 19705 18921 19717 18924
rect 19751 18921 19763 18955
rect 19705 18915 19763 18921
rect 22830 18912 22836 18964
rect 22888 18952 22894 18964
rect 25317 18955 25375 18961
rect 25317 18952 25329 18955
rect 22888 18924 25329 18952
rect 22888 18912 22894 18924
rect 25317 18921 25329 18924
rect 25363 18921 25375 18955
rect 25317 18915 25375 18921
rect 8938 18884 8944 18896
rect 8128 18856 8944 18884
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 3252 18816 3280 18856
rect 8938 18844 8944 18856
rect 8996 18844 9002 18896
rect 9030 18844 9036 18896
rect 9088 18884 9094 18896
rect 26053 18887 26111 18893
rect 26053 18884 26065 18887
rect 9088 18856 17172 18884
rect 9088 18844 9094 18856
rect 1903 18788 3280 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 3326 18776 3332 18828
rect 3384 18816 3390 18828
rect 14550 18816 14556 18828
rect 3384 18788 14556 18816
rect 3384 18776 3390 18788
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 15013 18819 15071 18825
rect 15013 18785 15025 18819
rect 15059 18816 15071 18819
rect 16758 18816 16764 18828
rect 15059 18788 16764 18816
rect 15059 18785 15071 18788
rect 15013 18779 15071 18785
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 1578 18748 1584 18760
rect 1539 18720 1584 18748
rect 1578 18708 1584 18720
rect 1636 18708 1642 18760
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 4157 18751 4215 18757
rect 4157 18748 4169 18751
rect 4028 18720 4169 18748
rect 4028 18708 4034 18720
rect 4157 18717 4169 18720
rect 4203 18717 4215 18751
rect 6546 18748 6552 18760
rect 5566 18720 6552 18748
rect 4157 18711 4215 18717
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 6822 18748 6828 18760
rect 6783 18720 6828 18748
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9953 18751 10011 18757
rect 9953 18717 9965 18751
rect 9999 18748 10011 18751
rect 10042 18748 10048 18760
rect 9999 18720 10048 18748
rect 9999 18717 10011 18720
rect 9953 18711 10011 18717
rect 3142 18680 3148 18692
rect 3082 18652 3148 18680
rect 3142 18640 3148 18652
rect 3200 18640 3206 18692
rect 4433 18683 4491 18689
rect 4433 18680 4445 18683
rect 3804 18652 4445 18680
rect 3804 18624 3832 18652
rect 4433 18649 4445 18652
rect 4479 18649 4491 18683
rect 7098 18680 7104 18692
rect 7059 18652 7104 18680
rect 4433 18643 4491 18649
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 7374 18640 7380 18692
rect 7432 18680 7438 18692
rect 7432 18652 7590 18680
rect 7432 18640 7438 18652
rect 3786 18572 3792 18624
rect 3844 18572 3850 18624
rect 5905 18615 5963 18621
rect 5905 18581 5917 18615
rect 5951 18612 5963 18615
rect 5994 18612 6000 18624
rect 5951 18584 6000 18612
rect 5951 18581 5963 18584
rect 5905 18575 5963 18581
rect 5994 18572 6000 18584
rect 6052 18572 6058 18624
rect 7466 18572 7472 18624
rect 7524 18612 7530 18624
rect 9324 18612 9352 18711
rect 10042 18708 10048 18720
rect 10100 18748 10106 18760
rect 10502 18748 10508 18760
rect 10100 18720 10508 18748
rect 10100 18708 10106 18720
rect 10502 18708 10508 18720
rect 10560 18708 10566 18760
rect 12158 18748 12164 18760
rect 12119 18720 12164 18748
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 12492 18720 13277 18748
rect 12492 18708 12498 18720
rect 13265 18717 13277 18720
rect 13311 18748 13323 18751
rect 14090 18748 14096 18760
rect 13311 18720 14096 18748
rect 13311 18717 13323 18720
rect 13265 18711 13323 18717
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18748 15531 18751
rect 16022 18748 16028 18760
rect 15519 18720 16028 18748
rect 15519 18717 15531 18720
rect 15473 18711 15531 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16390 18708 16396 18760
rect 16448 18748 16454 18760
rect 17144 18757 17172 18856
rect 25148 18856 26065 18884
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18816 23719 18819
rect 24026 18816 24032 18828
rect 23707 18788 24032 18816
rect 23707 18785 23719 18788
rect 23661 18779 23719 18785
rect 24026 18776 24032 18788
rect 24084 18776 24090 18828
rect 24946 18816 24952 18828
rect 24907 18788 24952 18816
rect 24946 18776 24952 18788
rect 25004 18776 25010 18828
rect 25148 18825 25176 18856
rect 26053 18853 26065 18856
rect 26099 18853 26111 18887
rect 38010 18884 38016 18896
rect 26053 18847 26111 18853
rect 31726 18856 38016 18884
rect 25133 18819 25191 18825
rect 25133 18785 25145 18819
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 16485 18751 16543 18757
rect 16485 18748 16497 18751
rect 16448 18720 16497 18748
rect 16448 18708 16454 18720
rect 16485 18717 16497 18720
rect 16531 18717 16543 18751
rect 16485 18711 16543 18717
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19978 18748 19984 18760
rect 19659 18720 19984 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20254 18748 20260 18760
rect 20215 18720 20260 18748
rect 20254 18708 20260 18720
rect 20312 18708 20318 18760
rect 25038 18708 25044 18760
rect 25096 18748 25102 18760
rect 26237 18751 26295 18757
rect 26237 18748 26249 18751
rect 25096 18720 26249 18748
rect 25096 18708 25102 18720
rect 26237 18717 26249 18720
rect 26283 18717 26295 18751
rect 26237 18711 26295 18717
rect 9582 18640 9588 18692
rect 9640 18680 9646 18692
rect 10686 18680 10692 18692
rect 9640 18652 10548 18680
rect 10647 18652 10692 18680
rect 9640 18640 9646 18652
rect 7524 18584 9352 18612
rect 7524 18572 7530 18584
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 10042 18612 10048 18624
rect 9456 18584 9501 18612
rect 10003 18584 10048 18612
rect 9456 18572 9462 18584
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10520 18612 10548 18652
rect 10686 18640 10692 18652
rect 10744 18640 10750 18692
rect 10778 18640 10784 18692
rect 10836 18680 10842 18692
rect 11698 18680 11704 18692
rect 10836 18652 10881 18680
rect 11659 18652 11704 18680
rect 10836 18640 10842 18652
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 13541 18683 13599 18689
rect 13541 18680 13553 18683
rect 12400 18652 13553 18680
rect 12400 18640 12406 18652
rect 13541 18649 13553 18652
rect 13587 18649 13599 18683
rect 13541 18643 13599 18649
rect 14182 18640 14188 18692
rect 14240 18680 14246 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 14240 18652 14381 18680
rect 14240 18640 14246 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 14461 18683 14519 18689
rect 14461 18649 14473 18683
rect 14507 18649 14519 18683
rect 14461 18643 14519 18649
rect 11974 18612 11980 18624
rect 10520 18584 11980 18612
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12253 18615 12311 18621
rect 12253 18581 12265 18615
rect 12299 18612 12311 18615
rect 14274 18612 14280 18624
rect 12299 18584 14280 18612
rect 12299 18581 12311 18584
rect 12253 18575 12311 18581
rect 14274 18572 14280 18584
rect 14332 18572 14338 18624
rect 14476 18612 14504 18643
rect 14550 18640 14556 18692
rect 14608 18680 14614 18692
rect 18414 18680 18420 18692
rect 14608 18652 18420 18680
rect 14608 18640 14614 18652
rect 18414 18640 18420 18652
rect 18472 18640 18478 18692
rect 22830 18640 22836 18692
rect 22888 18680 22894 18692
rect 23017 18683 23075 18689
rect 23017 18680 23029 18683
rect 22888 18652 23029 18680
rect 22888 18640 22894 18652
rect 23017 18649 23029 18652
rect 23063 18649 23075 18683
rect 23017 18643 23075 18649
rect 23109 18683 23167 18689
rect 23109 18649 23121 18683
rect 23155 18680 23167 18683
rect 23198 18680 23204 18692
rect 23155 18652 23204 18680
rect 23155 18649 23167 18652
rect 23109 18643 23167 18649
rect 23198 18640 23204 18652
rect 23256 18640 23262 18692
rect 31726 18680 31754 18856
rect 38010 18844 38016 18856
rect 38068 18844 38074 18896
rect 25516 18652 31754 18680
rect 16577 18615 16635 18621
rect 16577 18612 16589 18615
rect 14476 18584 16589 18612
rect 16577 18581 16589 18584
rect 16623 18581 16635 18615
rect 20346 18612 20352 18624
rect 20307 18584 20352 18612
rect 16577 18575 16635 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 20530 18572 20536 18624
rect 20588 18612 20594 18624
rect 25516 18612 25544 18652
rect 20588 18584 25544 18612
rect 20588 18572 20594 18584
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 3326 18408 3332 18420
rect 2832 18380 3332 18408
rect 2832 18368 2838 18380
rect 3326 18368 3332 18380
rect 3384 18368 3390 18420
rect 4062 18408 4068 18420
rect 3896 18380 4068 18408
rect 3896 18340 3924 18380
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 6822 18408 6828 18420
rect 4632 18380 6828 18408
rect 4632 18352 4660 18380
rect 4614 18340 4620 18352
rect 3082 18312 3924 18340
rect 4080 18312 4620 18340
rect 4080 18281 4108 18312
rect 4614 18300 4620 18312
rect 4672 18300 4678 18352
rect 4065 18275 4123 18281
rect 4065 18241 4077 18275
rect 4111 18241 4123 18275
rect 4065 18235 4123 18241
rect 5442 18232 5448 18284
rect 5500 18232 5506 18284
rect 6564 18281 6592 18380
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 8588 18380 11652 18408
rect 6730 18300 6736 18352
rect 6788 18340 6794 18352
rect 8588 18349 8616 18380
rect 8573 18343 8631 18349
rect 6788 18312 7314 18340
rect 6788 18300 6794 18312
rect 8573 18309 8585 18343
rect 8619 18309 8631 18343
rect 9306 18340 9312 18352
rect 9267 18312 9312 18340
rect 8573 18303 8631 18309
rect 9306 18300 9312 18312
rect 9364 18300 9370 18352
rect 10042 18300 10048 18352
rect 10100 18300 10106 18352
rect 11054 18300 11060 18352
rect 11112 18340 11118 18352
rect 11514 18340 11520 18352
rect 11112 18312 11520 18340
rect 11112 18300 11118 18312
rect 11514 18300 11520 18312
rect 11572 18300 11578 18352
rect 11624 18340 11652 18380
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 12986 18408 12992 18420
rect 11756 18380 12992 18408
rect 11756 18368 11762 18380
rect 12986 18368 12992 18380
rect 13044 18368 13050 18420
rect 14918 18408 14924 18420
rect 13096 18380 14924 18408
rect 11882 18340 11888 18352
rect 11624 18312 11888 18340
rect 11882 18300 11888 18312
rect 11940 18300 11946 18352
rect 11977 18343 12035 18349
rect 11977 18309 11989 18343
rect 12023 18340 12035 18343
rect 12066 18340 12072 18352
rect 12023 18312 12072 18340
rect 12023 18309 12035 18312
rect 11977 18303 12035 18309
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18241 6607 18275
rect 9033 18275 9091 18281
rect 9033 18272 9045 18275
rect 6549 18235 6607 18241
rect 8404 18244 9045 18272
rect 1578 18204 1584 18216
rect 1539 18176 1584 18204
rect 1578 18164 1584 18176
rect 1636 18164 1642 18216
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 3418 18204 3424 18216
rect 1903 18176 3424 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 4341 18207 4399 18213
rect 4341 18173 4353 18207
rect 4387 18204 4399 18207
rect 5718 18204 5724 18216
rect 4387 18176 5724 18204
rect 4387 18173 4399 18176
rect 4341 18167 4399 18173
rect 5718 18164 5724 18176
rect 5776 18164 5782 18216
rect 5813 18207 5871 18213
rect 5813 18173 5825 18207
rect 5859 18204 5871 18207
rect 6086 18204 6092 18216
rect 5859 18176 6092 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 6086 18164 6092 18176
rect 6144 18164 6150 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6196 18176 6837 18204
rect 2866 18096 2872 18148
rect 2924 18136 2930 18148
rect 6196 18136 6224 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 8404 18204 8432 18244
rect 6972 18176 8432 18204
rect 6972 18164 6978 18176
rect 2924 18108 4200 18136
rect 2924 18096 2930 18108
rect 4172 18068 4200 18108
rect 5368 18108 6224 18136
rect 8864 18136 8892 18244
rect 9033 18241 9045 18244
rect 9079 18241 9091 18275
rect 10778 18272 10784 18284
rect 9033 18235 9091 18241
rect 10520 18244 10784 18272
rect 8938 18164 8944 18216
rect 8996 18204 9002 18216
rect 9858 18204 9864 18216
rect 8996 18176 9864 18204
rect 8996 18164 9002 18176
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 9950 18164 9956 18216
rect 10008 18204 10014 18216
rect 10520 18204 10548 18244
rect 10778 18232 10784 18244
rect 10836 18232 10842 18284
rect 13096 18258 13124 18380
rect 14918 18368 14924 18380
rect 14976 18368 14982 18420
rect 15010 18368 15016 18420
rect 15068 18408 15074 18420
rect 21174 18408 21180 18420
rect 15068 18380 21180 18408
rect 15068 18368 15074 18380
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 23198 18408 23204 18420
rect 23159 18380 23204 18408
rect 23198 18368 23204 18380
rect 23256 18368 23262 18420
rect 23845 18411 23903 18417
rect 23845 18377 23857 18411
rect 23891 18408 23903 18411
rect 24394 18408 24400 18420
rect 23891 18380 24400 18408
rect 23891 18377 23903 18380
rect 23845 18371 23903 18377
rect 24394 18368 24400 18380
rect 24452 18368 24458 18420
rect 25038 18408 25044 18420
rect 24999 18380 25044 18408
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 14185 18343 14243 18349
rect 14185 18340 14197 18343
rect 13504 18312 14197 18340
rect 13504 18300 13510 18312
rect 14185 18309 14197 18312
rect 14231 18309 14243 18343
rect 14185 18303 14243 18309
rect 14274 18300 14280 18352
rect 14332 18340 14338 18352
rect 14332 18312 15700 18340
rect 14332 18300 14338 18312
rect 15010 18232 15016 18284
rect 15068 18232 15074 18284
rect 15672 18272 15700 18312
rect 18230 18300 18236 18352
rect 18288 18340 18294 18352
rect 19061 18343 19119 18349
rect 19061 18340 19073 18343
rect 18288 18312 19073 18340
rect 18288 18300 18294 18312
rect 19061 18309 19073 18312
rect 19107 18309 19119 18343
rect 19061 18303 19119 18309
rect 19153 18343 19211 18349
rect 19153 18309 19165 18343
rect 19199 18340 19211 18343
rect 20622 18340 20628 18352
rect 19199 18312 20628 18340
rect 19199 18309 19211 18312
rect 19153 18303 19211 18309
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15672 18244 15761 18272
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18049 18275 18107 18281
rect 18049 18272 18061 18275
rect 18012 18244 18061 18272
rect 18012 18232 18018 18244
rect 18049 18241 18061 18244
rect 18095 18241 18107 18275
rect 23382 18272 23388 18284
rect 23343 18244 23388 18272
rect 18049 18235 18107 18241
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 24026 18272 24032 18284
rect 23987 18244 24032 18272
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 25225 18275 25283 18281
rect 25225 18241 25237 18275
rect 25271 18241 25283 18275
rect 25682 18272 25688 18284
rect 25643 18244 25688 18272
rect 25225 18235 25283 18241
rect 10008 18176 10548 18204
rect 10008 18164 10014 18176
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11572 18176 11713 18204
rect 11572 18164 11578 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 11701 18167 11759 18173
rect 11808 18176 14105 18204
rect 10704 18136 10732 18164
rect 11808 18136 11836 18176
rect 14093 18173 14105 18176
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 14458 18164 14464 18216
rect 14516 18204 14522 18216
rect 15028 18204 15056 18232
rect 15105 18207 15163 18213
rect 15105 18204 15117 18207
rect 14516 18176 15117 18204
rect 14516 18164 14522 18176
rect 15105 18173 15117 18176
rect 15151 18173 15163 18207
rect 15105 18167 15163 18173
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 16942 18204 16948 18216
rect 15611 18176 16948 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 19242 18164 19248 18216
rect 19300 18204 19306 18216
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 19300 18176 19349 18204
rect 19300 18164 19306 18176
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 23566 18204 23572 18216
rect 21968 18176 23572 18204
rect 21968 18164 21974 18176
rect 23566 18164 23572 18176
rect 23624 18204 23630 18216
rect 25240 18204 25268 18235
rect 25682 18232 25688 18244
rect 25740 18232 25746 18284
rect 34422 18232 34428 18284
rect 34480 18272 34486 18284
rect 35345 18275 35403 18281
rect 35345 18272 35357 18275
rect 34480 18244 35357 18272
rect 34480 18232 34486 18244
rect 35345 18241 35357 18244
rect 35391 18241 35403 18275
rect 35345 18235 35403 18241
rect 35434 18232 35440 18284
rect 35492 18272 35498 18284
rect 38013 18275 38071 18281
rect 38013 18272 38025 18275
rect 35492 18244 38025 18272
rect 35492 18232 35498 18244
rect 38013 18241 38025 18244
rect 38059 18241 38071 18275
rect 38013 18235 38071 18241
rect 23624 18176 25268 18204
rect 23624 18164 23630 18176
rect 8864 18108 9168 18136
rect 10704 18108 11836 18136
rect 5368 18068 5396 18108
rect 4172 18040 5396 18068
rect 9140 18068 9168 18108
rect 15010 18096 15016 18148
rect 15068 18136 15074 18148
rect 19978 18136 19984 18148
rect 15068 18108 19984 18136
rect 15068 18096 15074 18108
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 10686 18068 10692 18080
rect 9140 18040 10692 18068
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 10781 18071 10839 18077
rect 10781 18037 10793 18071
rect 10827 18068 10839 18071
rect 10870 18068 10876 18080
rect 10827 18040 10876 18068
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 13446 18068 13452 18080
rect 11296 18040 13452 18068
rect 11296 18028 11302 18040
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 15930 18068 15936 18080
rect 13596 18040 15936 18068
rect 13596 18028 13602 18040
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16206 18068 16212 18080
rect 16167 18040 16212 18068
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 18141 18071 18199 18077
rect 18141 18037 18153 18071
rect 18187 18068 18199 18071
rect 18322 18068 18328 18080
rect 18187 18040 18328 18068
rect 18187 18037 18199 18040
rect 18141 18031 18199 18037
rect 18322 18028 18328 18040
rect 18380 18028 18386 18080
rect 25774 18068 25780 18080
rect 25735 18040 25780 18068
rect 25774 18028 25780 18040
rect 25832 18028 25838 18080
rect 35161 18071 35219 18077
rect 35161 18037 35173 18071
rect 35207 18068 35219 18071
rect 38010 18068 38016 18080
rect 35207 18040 38016 18068
rect 35207 18037 35219 18040
rect 35161 18031 35219 18037
rect 38010 18028 38016 18040
rect 38068 18028 38074 18080
rect 38194 18068 38200 18080
rect 38155 18040 38200 18068
rect 38194 18028 38200 18040
rect 38252 18028 38258 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 3970 17824 3976 17876
rect 4028 17824 4034 17876
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4120 17836 10732 17864
rect 4120 17824 4126 17836
rect 3050 17756 3056 17808
rect 3108 17796 3114 17808
rect 3421 17799 3479 17805
rect 3421 17796 3433 17799
rect 3108 17768 3433 17796
rect 3108 17756 3114 17768
rect 3421 17765 3433 17768
rect 3467 17796 3479 17799
rect 3786 17796 3792 17808
rect 3467 17768 3792 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 3988 17796 4016 17824
rect 3988 17768 4108 17796
rect 1670 17728 1676 17740
rect 1583 17700 1676 17728
rect 1670 17688 1676 17700
rect 1728 17728 1734 17740
rect 4080 17737 4108 17768
rect 5442 17756 5448 17808
rect 5500 17796 5506 17808
rect 10704 17796 10732 17836
rect 10778 17824 10784 17876
rect 10836 17864 10842 17876
rect 12066 17864 12072 17876
rect 10836 17836 12072 17864
rect 10836 17824 10842 17836
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 15838 17864 15844 17876
rect 12308 17836 15844 17864
rect 12308 17824 12314 17836
rect 15838 17824 15844 17836
rect 15896 17824 15902 17876
rect 15933 17867 15991 17873
rect 15933 17833 15945 17867
rect 15979 17864 15991 17867
rect 16574 17864 16580 17876
rect 15979 17836 16580 17864
rect 15979 17833 15991 17836
rect 15933 17827 15991 17833
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 18782 17864 18788 17876
rect 16684 17836 18788 17864
rect 16684 17796 16712 17836
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 22646 17796 22652 17808
rect 5500 17768 6960 17796
rect 10704 17768 11744 17796
rect 5500 17756 5506 17768
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 1728 17700 4077 17728
rect 1728 17688 1734 17700
rect 4065 17697 4077 17700
rect 4111 17728 4123 17731
rect 4706 17728 4712 17740
rect 4111 17700 4712 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 6822 17728 6828 17740
rect 6783 17700 6828 17728
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 6932 17728 6960 17768
rect 8573 17731 8631 17737
rect 8573 17728 8585 17731
rect 6932 17700 8585 17728
rect 8573 17697 8585 17700
rect 8619 17728 8631 17731
rect 8938 17728 8944 17740
rect 8619 17700 8944 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9125 17731 9183 17737
rect 9125 17697 9137 17731
rect 9171 17728 9183 17731
rect 11514 17728 11520 17740
rect 9171 17700 11520 17728
rect 9171 17697 9183 17700
rect 9125 17691 9183 17697
rect 11514 17688 11520 17700
rect 11572 17728 11578 17740
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11572 17700 11621 17728
rect 11572 17688 11578 17700
rect 11609 17697 11621 17700
rect 11655 17697 11667 17731
rect 11716 17728 11744 17768
rect 14384 17768 16712 17796
rect 17144 17768 22652 17796
rect 12250 17728 12256 17740
rect 11716 17700 12256 17728
rect 11609 17691 11667 17697
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 12342 17688 12348 17740
rect 12400 17728 12406 17740
rect 14384 17737 14412 17768
rect 13357 17731 13415 17737
rect 13357 17728 13369 17731
rect 12400 17700 13369 17728
rect 12400 17688 12406 17700
rect 13357 17697 13369 17700
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 14369 17731 14427 17737
rect 14369 17697 14381 17731
rect 14415 17697 14427 17731
rect 14369 17691 14427 17697
rect 15010 17688 15016 17740
rect 15068 17728 15074 17740
rect 15068 17700 16528 17728
rect 15068 17688 15074 17700
rect 10534 17632 11652 17660
rect 1946 17592 1952 17604
rect 1907 17564 1952 17592
rect 1946 17552 1952 17564
rect 2004 17552 2010 17604
rect 3174 17564 3832 17592
rect 3804 17524 3832 17564
rect 4246 17552 4252 17604
rect 4304 17592 4310 17604
rect 4341 17595 4399 17601
rect 4341 17592 4353 17595
rect 4304 17564 4353 17592
rect 4304 17552 4310 17564
rect 4341 17561 4353 17564
rect 4387 17561 4399 17595
rect 4341 17555 4399 17561
rect 5074 17552 5080 17604
rect 5132 17552 5138 17604
rect 7101 17595 7159 17601
rect 7101 17561 7113 17595
rect 7147 17561 7159 17595
rect 9306 17592 9312 17604
rect 8326 17564 9312 17592
rect 7101 17555 7159 17561
rect 4982 17524 4988 17536
rect 3804 17496 4988 17524
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 5813 17527 5871 17533
rect 5813 17493 5825 17527
rect 5859 17524 5871 17527
rect 5902 17524 5908 17536
rect 5859 17496 5908 17524
rect 5859 17493 5871 17496
rect 5813 17487 5871 17493
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 7116 17524 7144 17555
rect 9306 17552 9312 17564
rect 9364 17552 9370 17604
rect 9401 17595 9459 17601
rect 9401 17561 9413 17595
rect 9447 17561 9459 17595
rect 9401 17555 9459 17561
rect 9122 17524 9128 17536
rect 7116 17496 9128 17524
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 9416 17524 9444 17555
rect 10962 17552 10968 17604
rect 11020 17592 11026 17604
rect 11149 17595 11207 17601
rect 11149 17592 11161 17595
rect 11020 17564 11161 17592
rect 11020 17552 11026 17564
rect 11149 17561 11161 17564
rect 11195 17561 11207 17595
rect 11149 17555 11207 17561
rect 10870 17524 10876 17536
rect 9416 17496 10876 17524
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11624 17524 11652 17632
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 16500 17669 16528 17700
rect 17144 17669 17172 17768
rect 22646 17756 22652 17768
rect 22704 17756 22710 17808
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17728 19763 17731
rect 20346 17728 20352 17740
rect 19751 17700 20352 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 20346 17688 20352 17700
rect 20404 17728 20410 17740
rect 20809 17731 20867 17737
rect 20809 17728 20821 17731
rect 20404 17700 20821 17728
rect 20404 17688 20410 17700
rect 20809 17697 20821 17700
rect 20855 17697 20867 17731
rect 20809 17691 20867 17697
rect 20993 17731 21051 17737
rect 20993 17697 21005 17731
rect 21039 17728 21051 17731
rect 21266 17728 21272 17740
rect 21039 17700 21272 17728
rect 21039 17697 21051 17700
rect 20993 17691 21051 17697
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15344 17632 15853 17660
rect 15344 17620 15350 17632
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 11882 17552 11888 17604
rect 11940 17592 11946 17604
rect 13170 17592 13176 17604
rect 11940 17564 11985 17592
rect 13110 17564 13176 17592
rect 11940 17552 11946 17564
rect 13170 17552 13176 17564
rect 13228 17552 13234 17604
rect 14182 17592 14188 17604
rect 13740 17564 14188 17592
rect 13740 17524 13768 17564
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 14458 17552 14464 17604
rect 14516 17592 14522 17604
rect 15378 17592 15384 17604
rect 14516 17564 14561 17592
rect 15339 17564 15384 17592
rect 14516 17552 14522 17564
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 17494 17552 17500 17604
rect 17552 17592 17558 17604
rect 19797 17595 19855 17601
rect 17552 17564 19748 17592
rect 17552 17552 17558 17564
rect 11624 17496 13768 17524
rect 13814 17484 13820 17536
rect 13872 17524 13878 17536
rect 14826 17524 14832 17536
rect 13872 17496 14832 17524
rect 13872 17484 13878 17496
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 16574 17524 16580 17536
rect 16535 17496 16580 17524
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 17218 17524 17224 17536
rect 17179 17496 17224 17524
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 19720 17524 19748 17564
rect 19797 17561 19809 17595
rect 19843 17592 19855 17595
rect 20070 17592 20076 17604
rect 19843 17564 20076 17592
rect 19843 17561 19855 17564
rect 19797 17555 19855 17561
rect 20070 17552 20076 17564
rect 20128 17552 20134 17604
rect 20349 17595 20407 17601
rect 20349 17561 20361 17595
rect 20395 17561 20407 17595
rect 20349 17555 20407 17561
rect 20364 17524 20392 17555
rect 21450 17524 21456 17536
rect 19720 17496 20392 17524
rect 21411 17496 21456 17524
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 2590 17320 2596 17332
rect 1872 17292 2596 17320
rect 1872 17264 1900 17292
rect 2590 17280 2596 17292
rect 2648 17280 2654 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 4172 17292 6009 17320
rect 1854 17252 1860 17264
rect 1815 17224 1860 17252
rect 1854 17212 1860 17224
rect 1912 17212 1918 17264
rect 4062 17252 4068 17264
rect 3082 17224 4068 17252
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 3786 17184 3792 17196
rect 3528 17156 3792 17184
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 3528 17116 3556 17156
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 2004 17088 3556 17116
rect 2004 17076 2010 17088
rect 3602 17076 3608 17128
rect 3660 17116 3666 17128
rect 3660 17088 3705 17116
rect 3660 17076 3666 17088
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 3970 17048 3976 17060
rect 3016 17020 3976 17048
rect 3016 17008 3022 17020
rect 3970 17008 3976 17020
rect 4028 17008 4034 17060
rect 1486 16940 1492 16992
rect 1544 16980 1550 16992
rect 4172 16980 4200 17292
rect 5997 17289 6009 17292
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 6086 17280 6092 17332
rect 6144 17320 6150 17332
rect 6144 17292 9352 17320
rect 6144 17280 6150 17292
rect 4522 17252 4528 17264
rect 4483 17224 4528 17252
rect 4522 17212 4528 17224
rect 4580 17212 4586 17264
rect 9324 17252 9352 17292
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 10100 17292 14228 17320
rect 10100 17280 10106 17292
rect 9324 17224 10180 17252
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17116 4307 17119
rect 4614 17116 4620 17128
rect 4295 17088 4620 17116
rect 4295 17085 4307 17088
rect 4249 17079 4307 17085
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 4890 17076 4896 17128
rect 4948 17116 4954 17128
rect 6656 17116 6684 17147
rect 4948 17088 6684 17116
rect 4948 17076 4954 17088
rect 7098 17076 7104 17128
rect 7156 17116 7162 17128
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7156 17088 7757 17116
rect 7156 17076 7162 17088
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17116 8079 17119
rect 8570 17116 8576 17128
rect 8067 17088 8576 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 9140 17116 9168 17170
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 10042 17184 10048 17196
rect 9732 17156 10048 17184
rect 9732 17144 9738 17156
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 10152 17184 10180 17224
rect 10686 17212 10692 17264
rect 10744 17252 10750 17264
rect 10781 17255 10839 17261
rect 10781 17252 10793 17255
rect 10744 17224 10793 17252
rect 10744 17212 10750 17224
rect 10781 17221 10793 17224
rect 10827 17221 10839 17255
rect 11974 17252 11980 17264
rect 11935 17224 11980 17252
rect 10781 17215 10839 17221
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 12066 17212 12072 17264
rect 12124 17252 12130 17264
rect 14200 17261 14228 17292
rect 14458 17280 14464 17332
rect 14516 17320 14522 17332
rect 16945 17323 17003 17329
rect 16945 17320 16957 17323
rect 14516 17292 16957 17320
rect 14516 17280 14522 17292
rect 16945 17289 16957 17292
rect 16991 17289 17003 17323
rect 16945 17283 17003 17289
rect 34241 17323 34299 17329
rect 34241 17289 34253 17323
rect 34287 17320 34299 17323
rect 35434 17320 35440 17332
rect 34287 17292 35440 17320
rect 34287 17289 34299 17292
rect 34241 17283 34299 17289
rect 35434 17280 35440 17292
rect 35492 17280 35498 17332
rect 14185 17255 14243 17261
rect 12124 17224 12466 17252
rect 12124 17212 12130 17224
rect 14185 17221 14197 17255
rect 14231 17221 14243 17255
rect 14185 17215 14243 17221
rect 15194 17212 15200 17264
rect 15252 17252 15258 17264
rect 15657 17255 15715 17261
rect 15657 17252 15669 17255
rect 15252 17224 15669 17252
rect 15252 17212 15258 17224
rect 15657 17221 15669 17224
rect 15703 17221 15715 17255
rect 15657 17215 15715 17221
rect 15749 17255 15807 17261
rect 15749 17221 15761 17255
rect 15795 17252 15807 17255
rect 17218 17252 17224 17264
rect 15795 17224 17224 17252
rect 15795 17221 15807 17224
rect 15749 17215 15807 17221
rect 17218 17212 17224 17224
rect 17276 17212 17282 17264
rect 23109 17255 23167 17261
rect 23109 17221 23121 17255
rect 23155 17252 23167 17255
rect 23934 17252 23940 17264
rect 23155 17224 23940 17252
rect 23155 17221 23167 17224
rect 23109 17215 23167 17221
rect 23934 17212 23940 17224
rect 23992 17212 23998 17264
rect 24489 17255 24547 17261
rect 24489 17221 24501 17255
rect 24535 17252 24547 17255
rect 25774 17252 25780 17264
rect 24535 17224 25780 17252
rect 24535 17221 24547 17224
rect 24489 17215 24547 17221
rect 25774 17212 25780 17224
rect 25832 17212 25838 17264
rect 11330 17184 11336 17196
rect 10152 17156 11336 17184
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 10870 17116 10876 17128
rect 9140 17088 10876 17116
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 9306 17008 9312 17060
rect 9364 17048 9370 17060
rect 11606 17048 11612 17060
rect 9364 17020 11612 17048
rect 9364 17008 9370 17020
rect 11606 17008 11612 17020
rect 11664 17008 11670 17060
rect 1544 16952 4200 16980
rect 1544 16940 1550 16952
rect 5074 16940 5080 16992
rect 5132 16980 5138 16992
rect 6362 16980 6368 16992
rect 5132 16952 6368 16980
rect 5132 16940 5138 16952
rect 6362 16940 6368 16952
rect 6420 16940 6426 16992
rect 6730 16980 6736 16992
rect 6691 16952 6736 16980
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 11422 16980 11428 16992
rect 9539 16952 11428 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 11716 16980 11744 17147
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 16853 17187 16911 17193
rect 13688 17156 15056 17184
rect 13688 17144 13694 17156
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17116 13783 17119
rect 14734 17116 14740 17128
rect 13771 17088 14740 17116
rect 13771 17085 13783 17088
rect 13725 17079 13783 17085
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 14936 16980 14964 17079
rect 15028 17048 15056 17156
rect 16853 17153 16865 17187
rect 16899 17153 16911 17187
rect 17865 17187 17923 17193
rect 17865 17184 17877 17187
rect 16853 17147 16911 17153
rect 16960 17156 17877 17184
rect 16868 17116 16896 17147
rect 15764 17088 16896 17116
rect 15764 17048 15792 17088
rect 15028 17020 15792 17048
rect 16209 17051 16267 17057
rect 16209 17017 16221 17051
rect 16255 17017 16267 17051
rect 16209 17011 16267 17017
rect 11572 16952 14964 16980
rect 11572 16940 11578 16952
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 16224 16980 16252 17011
rect 16390 17008 16396 17060
rect 16448 17048 16454 17060
rect 16960 17048 16988 17156
rect 17865 17153 17877 17156
rect 17911 17153 17923 17187
rect 17865 17147 17923 17153
rect 19426 17144 19432 17196
rect 19484 17184 19490 17196
rect 20073 17187 20131 17193
rect 20073 17184 20085 17187
rect 19484 17156 20085 17184
rect 19484 17144 19490 17156
rect 20073 17153 20085 17156
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17184 23719 17187
rect 23750 17184 23756 17196
rect 23707 17156 23756 17184
rect 23707 17153 23719 17156
rect 23661 17147 23719 17153
rect 23750 17144 23756 17156
rect 23808 17144 23814 17196
rect 31754 17144 31760 17196
rect 31812 17184 31818 17196
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 31812 17156 34437 17184
rect 31812 17144 31818 17156
rect 34425 17153 34437 17156
rect 34471 17153 34483 17187
rect 34425 17147 34483 17153
rect 23014 17116 23020 17128
rect 22975 17088 23020 17116
rect 23014 17076 23020 17088
rect 23072 17076 23078 17128
rect 24394 17116 24400 17128
rect 24355 17088 24400 17116
rect 24394 17076 24400 17088
rect 24452 17076 24458 17128
rect 25409 17119 25467 17125
rect 25409 17085 25421 17119
rect 25455 17116 25467 17119
rect 25682 17116 25688 17128
rect 25455 17088 25688 17116
rect 25455 17085 25467 17088
rect 25409 17079 25467 17085
rect 25682 17076 25688 17088
rect 25740 17076 25746 17128
rect 16448 17020 16988 17048
rect 16448 17008 16454 17020
rect 17034 17008 17040 17060
rect 17092 17048 17098 17060
rect 24026 17048 24032 17060
rect 17092 17020 24032 17048
rect 17092 17008 17098 17020
rect 24026 17008 24032 17020
rect 24084 17008 24090 17060
rect 15436 16952 16252 16980
rect 15436 16940 15442 16952
rect 16850 16940 16856 16992
rect 16908 16980 16914 16992
rect 17678 16980 17684 16992
rect 16908 16952 17684 16980
rect 16908 16940 16914 16952
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 17957 16983 18015 16989
rect 17957 16949 17969 16983
rect 18003 16980 18015 16983
rect 18046 16980 18052 16992
rect 18003 16952 18052 16980
rect 18003 16949 18015 16952
rect 17957 16943 18015 16949
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 20162 16980 20168 16992
rect 20123 16952 20168 16980
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 26142 16980 26148 16992
rect 20956 16952 26148 16980
rect 20956 16940 20962 16952
rect 26142 16940 26148 16952
rect 26200 16940 26206 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1486 16736 1492 16788
rect 1544 16736 1550 16788
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 2038 16776 2044 16788
rect 1636 16748 2044 16776
rect 1636 16736 1642 16748
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 5708 16779 5766 16785
rect 5708 16745 5720 16779
rect 5754 16776 5766 16779
rect 6086 16776 6092 16788
rect 5754 16748 6092 16776
rect 5754 16745 5766 16748
rect 5708 16739 5766 16745
rect 6086 16736 6092 16748
rect 6144 16736 6150 16788
rect 6362 16736 6368 16788
rect 6420 16776 6426 16788
rect 6420 16748 9168 16776
rect 6420 16736 6426 16748
rect 1504 16708 1532 16736
rect 1504 16680 1808 16708
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 1780 16640 1808 16680
rect 4154 16668 4160 16720
rect 4212 16708 4218 16720
rect 4890 16708 4896 16720
rect 4212 16680 4896 16708
rect 4212 16668 4218 16680
rect 4890 16668 4896 16680
rect 4948 16668 4954 16720
rect 9140 16708 9168 16748
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 9364 16748 9409 16776
rect 9364 16736 9370 16748
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10597 16779 10655 16785
rect 10597 16776 10609 16779
rect 10008 16748 10609 16776
rect 10008 16736 10014 16748
rect 10597 16745 10609 16748
rect 10643 16745 10655 16779
rect 10597 16739 10655 16745
rect 11412 16779 11470 16785
rect 11412 16745 11424 16779
rect 11458 16776 11470 16779
rect 11790 16776 11796 16788
rect 11458 16748 11796 16776
rect 11458 16745 11470 16748
rect 11412 16739 11470 16745
rect 11790 16736 11796 16748
rect 11848 16776 11854 16788
rect 11848 16748 13124 16776
rect 11848 16736 11854 16748
rect 9140 16680 9536 16708
rect 1949 16643 2007 16649
rect 1949 16640 1961 16643
rect 1780 16612 1961 16640
rect 1949 16609 1961 16612
rect 1995 16609 2007 16643
rect 1949 16603 2007 16609
rect 3602 16600 3608 16652
rect 3660 16640 3666 16652
rect 3660 16612 4568 16640
rect 3660 16600 3666 16612
rect 3878 16572 3884 16584
rect 3082 16544 3884 16572
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4540 16572 4568 16612
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 5445 16643 5503 16649
rect 5445 16640 5457 16643
rect 4672 16612 5457 16640
rect 4672 16600 4678 16612
rect 5445 16609 5457 16612
rect 5491 16640 5503 16643
rect 7098 16640 7104 16652
rect 5491 16612 7104 16640
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 7098 16600 7104 16612
rect 7156 16640 7162 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 7156 16612 8401 16640
rect 7156 16600 7162 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 9508 16640 9536 16680
rect 9582 16668 9588 16720
rect 9640 16708 9646 16720
rect 11054 16708 11060 16720
rect 9640 16680 11060 16708
rect 9640 16668 9646 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 12710 16668 12716 16720
rect 12768 16708 12774 16720
rect 12894 16708 12900 16720
rect 12768 16680 12900 16708
rect 12768 16668 12774 16680
rect 12894 16668 12900 16680
rect 12952 16668 12958 16720
rect 13096 16708 13124 16748
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13228 16748 13645 16776
rect 13228 16736 13234 16748
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 13633 16739 13691 16745
rect 15838 16736 15844 16788
rect 15896 16776 15902 16788
rect 16025 16779 16083 16785
rect 16025 16776 16037 16779
rect 15896 16748 16037 16776
rect 15896 16736 15902 16748
rect 16025 16745 16037 16748
rect 16071 16745 16083 16779
rect 16025 16739 16083 16745
rect 16114 16736 16120 16788
rect 16172 16776 16178 16788
rect 19334 16776 19340 16788
rect 16172 16748 19340 16776
rect 16172 16736 16178 16748
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 37918 16776 37924 16788
rect 31726 16748 37924 16776
rect 17034 16708 17040 16720
rect 13096 16680 17040 16708
rect 17034 16668 17040 16680
rect 17092 16668 17098 16720
rect 31726 16708 31754 16748
rect 37918 16736 37924 16748
rect 37976 16736 37982 16788
rect 19812 16680 20116 16708
rect 11149 16643 11207 16649
rect 9508 16612 9904 16640
rect 8389 16603 8447 16609
rect 9209 16585 9267 16591
rect 5074 16572 5080 16584
rect 4540 16544 5080 16572
rect 5074 16532 5080 16544
rect 5132 16532 5138 16584
rect 8570 16532 8576 16584
rect 8628 16572 8634 16584
rect 9209 16582 9221 16585
rect 8956 16572 9221 16582
rect 8628 16554 9221 16572
rect 8628 16544 8984 16554
rect 9209 16551 9221 16554
rect 9255 16551 9267 16585
rect 9209 16545 9267 16551
rect 8628 16532 8634 16544
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 9876 16581 9904 16612
rect 11149 16609 11161 16643
rect 11195 16640 11207 16643
rect 11514 16640 11520 16652
rect 11195 16612 11520 16640
rect 11195 16609 11207 16612
rect 11149 16603 11207 16609
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 12158 16640 12164 16652
rect 11940 16612 12164 16640
rect 11940 16600 11946 16612
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 12986 16600 12992 16652
rect 13044 16640 13050 16652
rect 13354 16640 13360 16652
rect 13044 16612 13360 16640
rect 13044 16600 13050 16612
rect 13354 16600 13360 16612
rect 13412 16640 13418 16652
rect 16669 16643 16727 16649
rect 13412 16612 13492 16640
rect 13412 16600 13418 16612
rect 9861 16575 9919 16581
rect 9640 16532 9674 16572
rect 9861 16541 9873 16575
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10134 16572 10140 16584
rect 9999 16544 10140 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 10502 16532 10508 16584
rect 10560 16572 10566 16584
rect 10560 16544 10605 16572
rect 13464 16566 13492 16612
rect 16669 16609 16681 16643
rect 16715 16640 16727 16643
rect 16758 16640 16764 16652
rect 16715 16612 16764 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 18322 16640 18328 16652
rect 18283 16612 18328 16640
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 13541 16575 13599 16581
rect 13541 16566 13553 16575
rect 10560 16532 10566 16544
rect 13464 16541 13553 16566
rect 13587 16541 13599 16575
rect 13464 16538 13599 16541
rect 13541 16535 13599 16538
rect 14090 16532 14096 16584
rect 14148 16572 14154 16584
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14148 16544 14749 16572
rect 14148 16532 14154 16544
rect 14737 16541 14749 16544
rect 14783 16572 14795 16575
rect 14783 16544 15148 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 9646 16516 9674 16532
rect 3970 16504 3976 16516
rect 3931 16476 3976 16504
rect 3970 16464 3976 16476
rect 4028 16464 4034 16516
rect 4246 16464 4252 16516
rect 4304 16504 4310 16516
rect 4706 16504 4712 16516
rect 4304 16476 4712 16504
rect 4304 16464 4310 16476
rect 4706 16464 4712 16476
rect 4764 16464 4770 16516
rect 5626 16464 5632 16516
rect 5684 16504 5690 16516
rect 7650 16504 7656 16516
rect 5684 16476 6210 16504
rect 7024 16476 7656 16504
rect 5684 16464 5690 16476
rect 2866 16396 2872 16448
rect 2924 16436 2930 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 2924 16408 3433 16436
rect 2924 16396 2930 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3988 16436 4016 16464
rect 7024 16436 7052 16476
rect 7650 16464 7656 16476
rect 7708 16464 7714 16516
rect 9646 16476 9680 16516
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 11146 16504 11152 16516
rect 10428 16476 11152 16504
rect 3988 16408 7052 16436
rect 7193 16439 7251 16445
rect 3421 16399 3479 16405
rect 7193 16405 7205 16439
rect 7239 16436 7251 16439
rect 8018 16436 8024 16448
rect 7239 16408 8024 16436
rect 7239 16405 7251 16408
rect 7193 16399 7251 16405
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 10428 16436 10456 16476
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 14826 16504 14832 16516
rect 12650 16476 14832 16504
rect 14826 16464 14832 16476
rect 14884 16464 14890 16516
rect 15010 16504 15016 16516
rect 14971 16476 15016 16504
rect 15010 16464 15016 16476
rect 15068 16464 15074 16516
rect 15120 16504 15148 16544
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15933 16575 15991 16581
rect 15933 16572 15945 16575
rect 15620 16544 15945 16572
rect 15620 16532 15626 16544
rect 15933 16541 15945 16544
rect 15979 16541 15991 16575
rect 15933 16535 15991 16541
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16572 18199 16575
rect 18598 16572 18604 16584
rect 18187 16544 18604 16572
rect 18187 16541 18199 16544
rect 18141 16535 18199 16541
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 19812 16572 19840 16680
rect 18708 16544 19840 16572
rect 19889 16575 19947 16581
rect 15838 16504 15844 16516
rect 15120 16476 15844 16504
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 16758 16464 16764 16516
rect 16816 16504 16822 16516
rect 17678 16504 17684 16516
rect 16816 16476 16861 16504
rect 17639 16476 17684 16504
rect 16816 16464 16822 16476
rect 17678 16464 17684 16476
rect 17736 16464 17742 16516
rect 18708 16504 18736 16544
rect 19889 16541 19901 16575
rect 19935 16572 19947 16575
rect 19978 16572 19984 16584
rect 19935 16544 19984 16572
rect 19935 16541 19947 16544
rect 19889 16535 19947 16541
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 20088 16572 20116 16680
rect 23124 16680 31754 16708
rect 20640 16612 20944 16640
rect 20640 16572 20668 16612
rect 20806 16572 20812 16584
rect 20088 16544 20668 16572
rect 20767 16544 20812 16572
rect 20806 16532 20812 16544
rect 20864 16532 20870 16584
rect 20916 16572 20944 16612
rect 22186 16572 22192 16584
rect 20916 16544 22192 16572
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 22922 16532 22928 16584
rect 22980 16572 22986 16584
rect 23124 16581 23152 16680
rect 24026 16640 24032 16652
rect 23860 16612 24032 16640
rect 23860 16581 23888 16612
rect 24026 16600 24032 16612
rect 24084 16600 24090 16652
rect 24673 16643 24731 16649
rect 24673 16609 24685 16643
rect 24719 16640 24731 16643
rect 24854 16640 24860 16652
rect 24719 16612 24860 16640
rect 24719 16609 24731 16612
rect 24673 16603 24731 16609
rect 24854 16600 24860 16612
rect 24912 16640 24918 16652
rect 25498 16640 25504 16652
rect 24912 16612 25504 16640
rect 24912 16600 24918 16612
rect 25498 16600 25504 16612
rect 25556 16600 25562 16652
rect 26142 16640 26148 16652
rect 26103 16612 26148 16640
rect 26142 16600 26148 16612
rect 26200 16600 26206 16652
rect 26329 16643 26387 16649
rect 26329 16609 26341 16643
rect 26375 16640 26387 16643
rect 27706 16640 27712 16652
rect 26375 16612 27712 16640
rect 26375 16609 26387 16612
rect 26329 16603 26387 16609
rect 27706 16600 27712 16612
rect 27764 16600 27770 16652
rect 23109 16575 23167 16581
rect 23109 16572 23121 16575
rect 22980 16544 23121 16572
rect 22980 16532 22986 16544
rect 23109 16541 23121 16544
rect 23155 16541 23167 16575
rect 23109 16535 23167 16541
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16541 23903 16575
rect 23845 16535 23903 16541
rect 23934 16532 23940 16584
rect 23992 16572 23998 16584
rect 27801 16575 27859 16581
rect 27801 16572 27813 16575
rect 23992 16544 24037 16572
rect 26804 16544 27813 16572
rect 23992 16532 23998 16544
rect 17972 16476 18736 16504
rect 18785 16507 18843 16513
rect 17972 16448 18000 16476
rect 18785 16473 18797 16507
rect 18831 16504 18843 16507
rect 21450 16504 21456 16516
rect 18831 16476 21456 16504
rect 18831 16473 18843 16476
rect 18785 16467 18843 16473
rect 21450 16464 21456 16476
rect 21508 16464 21514 16516
rect 22204 16504 22232 16532
rect 23382 16504 23388 16516
rect 22204 16476 23388 16504
rect 23382 16464 23388 16476
rect 23440 16464 23446 16516
rect 24762 16464 24768 16516
rect 24820 16504 24826 16516
rect 25682 16504 25688 16516
rect 24820 16476 24865 16504
rect 25643 16476 25688 16504
rect 24820 16464 24826 16476
rect 25682 16464 25688 16476
rect 25740 16464 25746 16516
rect 26804 16448 26832 16544
rect 27801 16541 27813 16544
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 27893 16575 27951 16581
rect 27893 16541 27905 16575
rect 27939 16572 27951 16575
rect 31754 16572 31760 16584
rect 27939 16544 31760 16572
rect 27939 16541 27951 16544
rect 27893 16535 27951 16541
rect 31754 16532 31760 16544
rect 31812 16532 31818 16584
rect 38010 16572 38016 16584
rect 37971 16544 38016 16572
rect 38010 16532 38016 16544
rect 38068 16532 38074 16584
rect 9640 16408 10456 16436
rect 9640 16396 9646 16408
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 17954 16436 17960 16448
rect 10928 16408 17960 16436
rect 10928 16396 10934 16408
rect 17954 16396 17960 16408
rect 18012 16396 18018 16448
rect 19978 16436 19984 16448
rect 19939 16408 19984 16436
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 20254 16396 20260 16448
rect 20312 16436 20318 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20312 16408 20637 16436
rect 20312 16396 20318 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 20625 16399 20683 16405
rect 22002 16396 22008 16448
rect 22060 16436 22066 16448
rect 23201 16439 23259 16445
rect 23201 16436 23213 16439
rect 22060 16408 23213 16436
rect 22060 16396 22066 16408
rect 23201 16405 23213 16408
rect 23247 16436 23259 16439
rect 24394 16436 24400 16448
rect 23247 16408 24400 16436
rect 23247 16405 23259 16408
rect 23201 16399 23259 16405
rect 24394 16396 24400 16408
rect 24452 16396 24458 16448
rect 26786 16436 26792 16448
rect 26747 16408 26792 16436
rect 26786 16396 26792 16408
rect 26844 16396 26850 16448
rect 38194 16436 38200 16448
rect 38155 16408 38200 16436
rect 38194 16396 38200 16408
rect 38252 16396 38258 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 3513 16235 3571 16241
rect 3513 16201 3525 16235
rect 3559 16232 3571 16235
rect 3786 16232 3792 16244
rect 3559 16204 3792 16232
rect 3559 16201 3571 16204
rect 3513 16195 3571 16201
rect 3786 16192 3792 16204
rect 3844 16192 3850 16244
rect 5994 16232 6000 16244
rect 5907 16204 6000 16232
rect 5994 16192 6000 16204
rect 6052 16232 6058 16244
rect 9582 16232 9588 16244
rect 6052 16204 9588 16232
rect 6052 16192 6058 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 10778 16232 10784 16244
rect 10643 16204 10784 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 12894 16192 12900 16244
rect 12952 16232 12958 16244
rect 13262 16232 13268 16244
rect 12952 16204 13268 16232
rect 12952 16192 12958 16204
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 20806 16232 20812 16244
rect 14415 16204 19472 16232
rect 20767 16204 20812 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 3326 16164 3332 16176
rect 3266 16136 3332 16164
rect 3326 16124 3332 16136
rect 3384 16124 3390 16176
rect 5810 16164 5816 16176
rect 5750 16136 5816 16164
rect 5810 16124 5816 16136
rect 5868 16124 5874 16176
rect 7377 16167 7435 16173
rect 7377 16133 7389 16167
rect 7423 16164 7435 16167
rect 7650 16164 7656 16176
rect 7423 16136 7656 16164
rect 7423 16133 7435 16136
rect 7377 16127 7435 16133
rect 7650 16124 7656 16136
rect 7708 16124 7714 16176
rect 11330 16164 11336 16176
rect 8602 16136 11336 16164
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 12250 16164 12256 16176
rect 11440 16136 12256 16164
rect 1670 16056 1676 16108
rect 1728 16096 1734 16108
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 1728 16068 1777 16096
rect 1728 16056 1734 16068
rect 1765 16065 1777 16068
rect 1811 16065 1823 16099
rect 4246 16096 4252 16108
rect 4207 16068 4252 16096
rect 1765 16059 1823 16065
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 7098 16096 7104 16108
rect 7059 16068 7104 16096
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9766 16096 9772 16108
rect 9171 16068 9772 16096
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10410 16096 10416 16108
rect 9907 16068 10416 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 10410 16056 10416 16068
rect 10468 16056 10474 16108
rect 10502 16056 10508 16108
rect 10560 16096 10566 16108
rect 10560 16068 10605 16096
rect 10560 16056 10566 16068
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 16028 2099 16031
rect 2774 16028 2780 16040
rect 2087 16000 2780 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 5534 16028 5540 16040
rect 4571 16000 5540 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 6236 16000 9904 16028
rect 6236 15988 6242 16000
rect 9876 15972 9904 16000
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 11440 16028 11468 16136
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 13202 16136 13768 16164
rect 10376 16000 11468 16028
rect 10376 15988 10382 16000
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 11572 16000 11713 16028
rect 11572 15988 11578 16000
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 13354 16028 13360 16040
rect 12023 16000 13360 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 9858 15920 9864 15972
rect 9916 15920 9922 15972
rect 9953 15963 10011 15969
rect 9953 15929 9965 15963
rect 9999 15960 10011 15963
rect 9999 15932 11836 15960
rect 9999 15929 10011 15932
rect 9953 15923 10011 15929
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 9122 15892 9128 15904
rect 6144 15864 9128 15892
rect 6144 15852 6150 15864
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 9214 15852 9220 15904
rect 9272 15892 9278 15904
rect 10318 15892 10324 15904
rect 9272 15864 10324 15892
rect 9272 15852 9278 15864
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 11808 15892 11836 15932
rect 11974 15892 11980 15904
rect 11808 15864 11980 15892
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 13412 15864 13461 15892
rect 13412 15852 13418 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13740 15892 13768 16136
rect 14826 16124 14832 16176
rect 14884 16164 14890 16176
rect 15749 16167 15807 16173
rect 15749 16164 15761 16167
rect 14884 16136 15761 16164
rect 14884 16124 14890 16136
rect 15749 16133 15761 16136
rect 15795 16133 15807 16167
rect 15749 16127 15807 16133
rect 17037 16167 17095 16173
rect 17037 16133 17049 16167
rect 17083 16164 17095 16167
rect 17310 16164 17316 16176
rect 17083 16136 17316 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 19444 16173 19472 16204
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 24762 16192 24768 16244
rect 24820 16232 24826 16244
rect 26329 16235 26387 16241
rect 26329 16232 26341 16235
rect 24820 16204 26341 16232
rect 24820 16192 24826 16204
rect 26329 16201 26341 16204
rect 26375 16201 26387 16235
rect 27706 16232 27712 16244
rect 27667 16204 27712 16232
rect 26329 16195 26387 16201
rect 27706 16192 27712 16204
rect 27764 16192 27770 16244
rect 28261 16235 28319 16241
rect 28261 16201 28273 16235
rect 28307 16201 28319 16235
rect 28261 16195 28319 16201
rect 19429 16167 19487 16173
rect 19429 16133 19441 16167
rect 19475 16133 19487 16167
rect 22186 16164 22192 16176
rect 22147 16136 22192 16164
rect 19429 16127 19487 16133
rect 22186 16124 22192 16136
rect 22244 16124 22250 16176
rect 28276 16164 28304 16195
rect 28276 16136 29132 16164
rect 14274 16096 14280 16108
rect 14235 16068 14280 16096
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14792 16068 14933 16096
rect 14792 16056 14798 16068
rect 14921 16065 14933 16068
rect 14967 16096 14979 16099
rect 15562 16096 15568 16108
rect 14967 16068 15568 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 15838 16096 15844 16108
rect 15703 16068 15844 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15838 16056 15844 16068
rect 15896 16096 15902 16108
rect 16298 16096 16304 16108
rect 15896 16068 16304 16096
rect 15896 16056 15902 16068
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 18966 16096 18972 16108
rect 18432 16068 18972 16096
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 15013 16031 15071 16037
rect 15013 16028 15025 16031
rect 13872 16000 15025 16028
rect 13872 15988 13878 16000
rect 15013 15997 15025 16000
rect 15059 15997 15071 16031
rect 16574 16028 16580 16040
rect 15013 15991 15071 15997
rect 15304 16000 16580 16028
rect 14550 15920 14556 15972
rect 14608 15960 14614 15972
rect 15304 15960 15332 16000
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 18432 16028 18460 16068
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 20993 16099 21051 16105
rect 20993 16096 21005 16099
rect 20180 16068 21005 16096
rect 16991 16000 18460 16028
rect 18601 16031 18659 16037
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 18601 15997 18613 16031
rect 18647 16028 18659 16031
rect 19337 16031 19395 16037
rect 19337 16028 19349 16031
rect 18647 16000 19349 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 19337 15997 19349 16000
rect 19383 15997 19395 16031
rect 19337 15991 19395 15997
rect 19426 15988 19432 16040
rect 19484 16028 19490 16040
rect 20180 16028 20208 16068
rect 20993 16065 21005 16068
rect 21039 16065 21051 16099
rect 26234 16096 26240 16108
rect 26195 16068 26240 16096
rect 20993 16059 21051 16065
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 27614 16096 27620 16108
rect 27575 16068 27620 16096
rect 27614 16056 27620 16068
rect 27672 16096 27678 16108
rect 29104 16105 29132 16136
rect 28445 16099 28503 16105
rect 28445 16096 28457 16099
rect 27672 16068 28457 16096
rect 27672 16056 27678 16068
rect 28445 16065 28457 16068
rect 28491 16065 28503 16099
rect 28445 16059 28503 16065
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16065 29147 16099
rect 29089 16059 29147 16065
rect 36538 16056 36544 16108
rect 36596 16096 36602 16108
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 36596 16068 38025 16096
rect 36596 16056 36602 16068
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 19484 16000 20208 16028
rect 20257 16031 20315 16037
rect 19484 15988 19490 16000
rect 20257 15997 20269 16031
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 14608 15932 15332 15960
rect 14608 15920 14614 15932
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 17494 15960 17500 15972
rect 15436 15932 17500 15960
rect 15436 15920 15442 15932
rect 17494 15920 17500 15932
rect 17552 15920 17558 15972
rect 17678 15920 17684 15972
rect 17736 15960 17742 15972
rect 18874 15960 18880 15972
rect 17736 15932 18880 15960
rect 17736 15920 17742 15932
rect 18874 15920 18880 15932
rect 18932 15960 18938 15972
rect 20272 15960 20300 15991
rect 21818 15988 21824 16040
rect 21876 16028 21882 16040
rect 22097 16031 22155 16037
rect 22097 16028 22109 16031
rect 21876 16000 22109 16028
rect 21876 15988 21882 16000
rect 22097 15997 22109 16000
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 22373 16031 22431 16037
rect 22373 15997 22385 16031
rect 22419 15997 22431 16031
rect 22373 15991 22431 15997
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 16028 24271 16031
rect 24578 16028 24584 16040
rect 24259 16000 24584 16028
rect 24259 15997 24271 16000
rect 24213 15991 24271 15997
rect 18932 15932 20300 15960
rect 18932 15920 18938 15932
rect 21726 15920 21732 15972
rect 21784 15960 21790 15972
rect 22388 15960 22416 15991
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 25682 15960 25688 15972
rect 21784 15932 22416 15960
rect 24688 15932 25688 15960
rect 21784 15920 21790 15932
rect 18506 15892 18512 15904
rect 13740 15864 18512 15892
rect 13449 15855 13507 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 18690 15852 18696 15904
rect 18748 15892 18754 15904
rect 24688 15892 24716 15932
rect 25682 15920 25688 15932
rect 25740 15920 25746 15972
rect 18748 15864 24716 15892
rect 18748 15852 18754 15864
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 28905 15895 28963 15901
rect 28905 15892 28917 15895
rect 24820 15864 28917 15892
rect 24820 15852 24826 15864
rect 28905 15861 28917 15864
rect 28951 15861 28963 15895
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 28905 15855 28963 15861
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 3329 15691 3387 15697
rect 3329 15657 3341 15691
rect 3375 15688 3387 15691
rect 3602 15688 3608 15700
rect 3375 15660 3608 15688
rect 3375 15657 3387 15660
rect 3329 15651 3387 15657
rect 3602 15648 3608 15660
rect 3660 15648 3666 15700
rect 4236 15691 4294 15697
rect 4236 15657 4248 15691
rect 4282 15688 4294 15691
rect 7190 15688 7196 15700
rect 4282 15660 7196 15688
rect 4282 15657 4294 15660
rect 4236 15651 4294 15657
rect 7190 15648 7196 15660
rect 7248 15688 7254 15700
rect 11790 15688 11796 15700
rect 7248 15660 11652 15688
rect 11751 15660 11796 15688
rect 7248 15648 7254 15660
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 5721 15623 5779 15629
rect 5721 15620 5733 15623
rect 5592 15592 5733 15620
rect 5592 15580 5598 15592
rect 5721 15589 5733 15592
rect 5767 15620 5779 15623
rect 6086 15620 6092 15632
rect 5767 15592 6092 15620
rect 5767 15589 5779 15592
rect 5721 15583 5779 15589
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 11624 15620 11652 15660
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 14734 15688 14740 15700
rect 12492 15660 14740 15688
rect 12492 15648 12498 15660
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 16574 15648 16580 15700
rect 16632 15688 16638 15700
rect 21726 15688 21732 15700
rect 16632 15660 21732 15688
rect 16632 15648 16638 15660
rect 21726 15648 21732 15660
rect 21784 15648 21790 15700
rect 22462 15688 22468 15700
rect 22375 15660 22468 15688
rect 22462 15648 22468 15660
rect 22520 15688 22526 15700
rect 23014 15688 23020 15700
rect 22520 15660 23020 15688
rect 22520 15648 22526 15660
rect 23014 15648 23020 15660
rect 23072 15648 23078 15700
rect 25225 15691 25283 15697
rect 25225 15657 25237 15691
rect 25271 15688 25283 15691
rect 26786 15688 26792 15700
rect 25271 15660 26792 15688
rect 25271 15657 25283 15660
rect 25225 15651 25283 15657
rect 26786 15648 26792 15660
rect 26844 15648 26850 15700
rect 13538 15620 13544 15632
rect 11624 15592 13544 15620
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 15562 15620 15568 15632
rect 15523 15592 15568 15620
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 20806 15620 20812 15632
rect 19260 15592 20812 15620
rect 1578 15552 1584 15564
rect 1539 15524 1584 15552
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 3418 15552 3424 15564
rect 1903 15524 3424 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 4614 15552 4620 15564
rect 3988 15524 4620 15552
rect 3988 15493 4016 15524
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15552 6607 15555
rect 6822 15552 6828 15564
rect 6595 15524 6828 15552
rect 6595 15521 6607 15524
rect 6549 15515 6607 15521
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 10686 15552 10692 15564
rect 10091 15524 10692 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 11606 15512 11612 15564
rect 11664 15552 11670 15564
rect 12802 15552 12808 15564
rect 11664 15524 12808 15552
rect 11664 15512 11670 15524
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 13170 15512 13176 15564
rect 13228 15552 13234 15564
rect 18690 15552 18696 15564
rect 13228 15524 13584 15552
rect 13228 15512 13234 15524
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 3988 15416 4016 15447
rect 5350 15444 5356 15496
rect 5408 15444 5414 15496
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 4154 15416 4160 15428
rect 3082 15388 3924 15416
rect 3988 15388 4160 15416
rect 1946 15308 1952 15360
rect 2004 15348 2010 15360
rect 2590 15348 2596 15360
rect 2004 15320 2596 15348
rect 2004 15308 2010 15320
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 3896 15348 3924 15388
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 6454 15376 6460 15428
rect 6512 15416 6518 15428
rect 6730 15416 6736 15428
rect 6512 15388 6736 15416
rect 6512 15376 6518 15388
rect 6730 15376 6736 15388
rect 6788 15376 6794 15428
rect 6825 15419 6883 15425
rect 6825 15385 6837 15419
rect 6871 15385 6883 15419
rect 6825 15379 6883 15385
rect 6178 15348 6184 15360
rect 3896 15320 6184 15348
rect 6178 15308 6184 15320
rect 6236 15308 6242 15360
rect 6840 15348 6868 15379
rect 7834 15376 7840 15428
rect 7892 15376 7898 15428
rect 9416 15416 9444 15447
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12526 15484 12532 15496
rect 12308 15456 12532 15484
rect 12308 15444 12314 15456
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13556 15484 13584 15524
rect 14752 15524 18696 15552
rect 14752 15484 14780 15524
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 13556 15456 14780 15484
rect 14829 15487 14887 15493
rect 9416 15388 10272 15416
rect 6914 15348 6920 15360
rect 6827 15320 6920 15348
rect 6914 15308 6920 15320
rect 6972 15348 6978 15360
rect 7742 15348 7748 15360
rect 6972 15320 7748 15348
rect 6972 15308 6978 15320
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 8297 15351 8355 15357
rect 8297 15317 8309 15351
rect 8343 15348 8355 15351
rect 8478 15348 8484 15360
rect 8343 15320 8484 15348
rect 8343 15317 8355 15320
rect 8297 15311 8355 15317
rect 8478 15308 8484 15320
rect 8536 15308 8542 15360
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9582 15348 9588 15360
rect 9539 15320 9588 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 10244 15348 10272 15388
rect 10318 15376 10324 15428
rect 10376 15416 10382 15428
rect 10376 15388 10421 15416
rect 10376 15376 10382 15388
rect 11054 15376 11060 15428
rect 11112 15376 11118 15428
rect 12713 15419 12771 15425
rect 12713 15385 12725 15419
rect 12759 15385 12771 15419
rect 12713 15379 12771 15385
rect 12805 15419 12863 15425
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 12894 15416 12900 15428
rect 12851 15388 12900 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 12434 15348 12440 15360
rect 10244 15320 12440 15348
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 12728 15348 12756 15379
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 13556 15348 13584 15456
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 14875 15456 15148 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 13725 15419 13783 15425
rect 13725 15385 13737 15419
rect 13771 15416 13783 15419
rect 15010 15416 15016 15428
rect 13771 15388 15016 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 15010 15376 15016 15388
rect 15068 15376 15074 15428
rect 15120 15416 15148 15456
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15252 15456 15485 15484
rect 15252 15444 15258 15456
rect 15473 15453 15485 15456
rect 15519 15453 15531 15487
rect 16114 15484 16120 15496
rect 16075 15456 16120 15484
rect 15473 15447 15531 15453
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 15286 15416 15292 15428
rect 15120 15388 15292 15416
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 15838 15376 15844 15428
rect 15896 15416 15902 15428
rect 17236 15416 17264 15447
rect 17310 15444 17316 15496
rect 17368 15484 17374 15496
rect 17862 15484 17868 15496
rect 17368 15456 17413 15484
rect 17823 15456 17868 15484
rect 17368 15444 17374 15456
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18472 15456 18521 15484
rect 18472 15444 18478 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 19260 15416 19288 15592
rect 20806 15580 20812 15592
rect 20864 15620 20870 15632
rect 21542 15620 21548 15632
rect 20864 15592 21548 15620
rect 20864 15580 20870 15592
rect 21542 15580 21548 15592
rect 21600 15580 21606 15632
rect 22925 15623 22983 15629
rect 22925 15620 22937 15623
rect 22112 15592 22937 15620
rect 21818 15484 21824 15496
rect 21779 15456 21824 15484
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 22005 15487 22063 15493
rect 22005 15453 22017 15487
rect 22051 15484 22063 15487
rect 22112 15484 22140 15592
rect 22925 15589 22937 15592
rect 22971 15589 22983 15623
rect 22925 15583 22983 15589
rect 23382 15580 23388 15632
rect 23440 15620 23446 15632
rect 27982 15620 27988 15632
rect 23440 15592 27988 15620
rect 23440 15580 23446 15592
rect 27982 15580 27988 15592
rect 28040 15620 28046 15632
rect 28040 15592 28764 15620
rect 28040 15580 28046 15592
rect 24578 15552 24584 15564
rect 22051 15456 22140 15484
rect 23032 15524 23796 15552
rect 24539 15524 24584 15552
rect 22051 15453 22063 15456
rect 22005 15447 22063 15453
rect 15896 15388 17264 15416
rect 17788 15388 19288 15416
rect 15896 15376 15902 15388
rect 12728 15320 13584 15348
rect 14826 15308 14832 15360
rect 14884 15348 14890 15360
rect 14921 15351 14979 15357
rect 14921 15348 14933 15351
rect 14884 15320 14933 15348
rect 14884 15308 14890 15320
rect 14921 15317 14933 15320
rect 14967 15317 14979 15351
rect 14921 15311 14979 15317
rect 16209 15351 16267 15357
rect 16209 15317 16221 15351
rect 16255 15348 16267 15351
rect 17034 15348 17040 15360
rect 16255 15320 17040 15348
rect 16255 15317 16267 15320
rect 16209 15311 16267 15317
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17126 15308 17132 15360
rect 17184 15348 17190 15360
rect 17788 15348 17816 15388
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19521 15419 19579 15425
rect 19521 15416 19533 15419
rect 19392 15388 19533 15416
rect 19392 15376 19398 15388
rect 19521 15385 19533 15388
rect 19567 15385 19579 15419
rect 19521 15379 19579 15385
rect 19613 15419 19671 15425
rect 19613 15385 19625 15419
rect 19659 15416 19671 15419
rect 19978 15416 19984 15428
rect 19659 15388 19984 15416
rect 19659 15385 19671 15388
rect 19613 15379 19671 15385
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 20165 15419 20223 15425
rect 20165 15385 20177 15419
rect 20211 15416 20223 15419
rect 20346 15416 20352 15428
rect 20211 15388 20352 15416
rect 20211 15385 20223 15388
rect 20165 15379 20223 15385
rect 20346 15376 20352 15388
rect 20404 15376 20410 15428
rect 21177 15419 21235 15425
rect 21177 15385 21189 15419
rect 21223 15416 21235 15419
rect 22922 15416 22928 15428
rect 21223 15388 22928 15416
rect 21223 15385 21235 15388
rect 21177 15379 21235 15385
rect 22922 15376 22928 15388
rect 22980 15376 22986 15428
rect 17954 15348 17960 15360
rect 17184 15320 17816 15348
rect 17915 15320 17960 15348
rect 17184 15308 17190 15320
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 18598 15348 18604 15360
rect 18559 15320 18604 15348
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 23032 15348 23060 15524
rect 23768 15493 23796 15524
rect 24578 15512 24584 15524
rect 24636 15512 24642 15564
rect 24762 15552 24768 15564
rect 24723 15524 24768 15552
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 28736 15493 28764 15592
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15484 23167 15487
rect 23753 15487 23811 15493
rect 23155 15456 23612 15484
rect 23155 15453 23167 15456
rect 23109 15447 23167 15453
rect 23584 15357 23612 15456
rect 23753 15453 23765 15487
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 28721 15487 28779 15493
rect 28721 15453 28733 15487
rect 28767 15453 28779 15487
rect 28721 15447 28779 15453
rect 21600 15320 23060 15348
rect 23569 15351 23627 15357
rect 21600 15308 21606 15320
rect 23569 15317 23581 15351
rect 23615 15317 23627 15351
rect 23569 15311 23627 15317
rect 28537 15351 28595 15357
rect 28537 15317 28549 15351
rect 28583 15348 28595 15351
rect 28810 15348 28816 15360
rect 28583 15320 28816 15348
rect 28583 15317 28595 15320
rect 28537 15311 28595 15317
rect 28810 15308 28816 15320
rect 28868 15308 28874 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 3602 15144 3608 15156
rect 1872 15116 3608 15144
rect 1872 15085 1900 15116
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 8478 15144 8484 15156
rect 4264 15116 8484 15144
rect 1857 15079 1915 15085
rect 1857 15045 1869 15079
rect 1903 15045 1915 15079
rect 4154 15076 4160 15088
rect 1857 15039 1915 15045
rect 3988 15048 4160 15076
rect 1578 15008 1584 15020
rect 1539 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 3988 15017 4016 15048
rect 4154 15036 4160 15048
rect 4212 15036 4218 15088
rect 4264 15085 4292 15116
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 9122 15104 9128 15156
rect 9180 15144 9186 15156
rect 9180 15116 9674 15144
rect 9180 15104 9186 15116
rect 4249 15079 4307 15085
rect 4249 15045 4261 15079
rect 4295 15045 4307 15079
rect 4249 15039 4307 15045
rect 4982 15036 4988 15088
rect 5040 15036 5046 15088
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 7892 15048 8786 15076
rect 7892 15036 7898 15048
rect 3973 15011 4031 15017
rect 2406 14900 2412 14952
rect 2464 14940 2470 14952
rect 2590 14940 2596 14952
rect 2464 14912 2596 14940
rect 2464 14900 2470 14912
rect 2590 14900 2596 14912
rect 2648 14900 2654 14952
rect 2976 14872 3004 14994
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7098 15008 7104 15020
rect 6963 14980 7104 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7466 15008 7472 15020
rect 7423 14980 7472 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 9646 15008 9674 15116
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 11057 15147 11115 15153
rect 10008 15116 11008 15144
rect 10008 15104 10014 15116
rect 10045 15079 10103 15085
rect 10045 15045 10057 15079
rect 10091 15076 10103 15079
rect 10226 15076 10232 15088
rect 10091 15048 10232 15076
rect 10091 15045 10103 15048
rect 10045 15039 10103 15045
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 10980 15076 11008 15116
rect 11057 15113 11069 15147
rect 11103 15144 11115 15147
rect 12894 15144 12900 15156
rect 11103 15116 12900 15144
rect 11103 15113 11115 15116
rect 11057 15107 11115 15113
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13412 15116 13461 15144
rect 13412 15104 13418 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 17954 15144 17960 15156
rect 13449 15107 13507 15113
rect 14200 15116 17960 15144
rect 14200 15085 14228 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18506 15144 18512 15156
rect 18467 15116 18512 15144
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 20714 15144 20720 15156
rect 20675 15116 20720 15144
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 22097 15147 22155 15153
rect 22097 15113 22109 15147
rect 22143 15144 22155 15147
rect 22186 15144 22192 15156
rect 22143 15116 22192 15144
rect 22143 15113 22155 15116
rect 22097 15107 22155 15113
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 14185 15079 14243 15085
rect 10980 15048 12466 15076
rect 14185 15045 14197 15079
rect 14231 15045 14243 15079
rect 14185 15039 14243 15045
rect 15010 15036 15016 15088
rect 15068 15076 15074 15088
rect 15105 15079 15163 15085
rect 15105 15076 15117 15079
rect 15068 15048 15117 15076
rect 15068 15036 15074 15048
rect 15105 15045 15117 15048
rect 15151 15045 15163 15079
rect 17034 15076 17040 15088
rect 16995 15048 17040 15076
rect 15105 15039 15163 15045
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20898 15076 20904 15088
rect 19935 15048 20904 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 21818 15036 21824 15088
rect 21876 15076 21882 15088
rect 24121 15079 24179 15085
rect 24121 15076 24133 15079
rect 21876 15048 24133 15076
rect 21876 15036 21882 15048
rect 24121 15045 24133 15048
rect 24167 15045 24179 15079
rect 24121 15039 24179 15045
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 9646 14980 10977 15008
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 18414 15008 18420 15020
rect 18375 14980 18420 15008
rect 10965 14971 11023 14977
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 15008 19487 15011
rect 20162 15008 20168 15020
rect 19475 14980 20168 15008
rect 19475 14977 19487 14980
rect 19429 14971 19487 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 15008 20683 15011
rect 21266 15008 21272 15020
rect 20671 14980 21272 15008
rect 20671 14977 20683 14980
rect 20625 14971 20683 14977
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 22002 15008 22008 15020
rect 21963 14980 22008 15008
rect 22002 14968 22008 14980
rect 22060 14968 22066 15020
rect 23842 14968 23848 15020
rect 23900 15008 23906 15020
rect 24029 15011 24087 15017
rect 24029 15008 24041 15011
rect 23900 14980 24041 15008
rect 23900 14968 23906 14980
rect 24029 14977 24041 14980
rect 24075 15008 24087 15011
rect 26050 15008 26056 15020
rect 24075 14980 26056 15008
rect 24075 14977 24087 14980
rect 24029 14971 24087 14977
rect 26050 14968 26056 14980
rect 26108 14968 26114 15020
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 26160 14980 26249 15008
rect 26160 14952 26188 14980
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 28810 15008 28816 15020
rect 28771 14980 28816 15008
rect 26237 14971 26295 14977
rect 28810 14968 28816 14980
rect 28868 14968 28874 15020
rect 37826 14968 37832 15020
rect 37884 15008 37890 15020
rect 38013 15011 38071 15017
rect 38013 15008 38025 15011
rect 37884 14980 38025 15008
rect 37884 14968 37890 14980
rect 38013 14977 38025 14980
rect 38059 14977 38071 15011
rect 38013 14971 38071 14977
rect 3326 14940 3332 14952
rect 3287 14912 3332 14940
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 5718 14940 5724 14952
rect 5679 14912 5724 14940
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 8021 14943 8079 14949
rect 8021 14940 8033 14943
rect 6880 14912 8033 14940
rect 6880 14900 6886 14912
rect 8021 14909 8033 14912
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 8297 14943 8355 14949
rect 8297 14909 8309 14943
rect 8343 14940 8355 14943
rect 9950 14940 9956 14952
rect 8343 14912 9956 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 11572 14912 11713 14940
rect 11572 14900 11578 14912
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12066 14940 12072 14952
rect 12023 14912 12072 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 15562 14940 15568 14952
rect 14139 14912 15568 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14940 16175 14943
rect 16945 14943 17003 14949
rect 16945 14940 16957 14943
rect 16163 14912 16957 14940
rect 16163 14909 16175 14912
rect 16117 14903 16175 14909
rect 16945 14909 16957 14912
rect 16991 14909 17003 14943
rect 17586 14940 17592 14952
rect 17547 14912 17592 14940
rect 16945 14903 17003 14909
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14940 19303 14943
rect 19334 14940 19340 14952
rect 19291 14912 19340 14940
rect 19291 14909 19303 14912
rect 19245 14903 19303 14909
rect 19334 14900 19340 14912
rect 19392 14940 19398 14952
rect 21361 14943 21419 14949
rect 21361 14940 21373 14943
rect 19392 14912 21373 14940
rect 19392 14900 19398 14912
rect 21361 14909 21373 14912
rect 21407 14909 21419 14943
rect 26142 14940 26148 14952
rect 21361 14903 21419 14909
rect 22066 14912 26148 14940
rect 6733 14875 6791 14881
rect 2976 14844 4016 14872
rect 3988 14804 4016 14844
rect 6733 14841 6745 14875
rect 6779 14872 6791 14875
rect 7006 14872 7012 14884
rect 6779 14844 7012 14872
rect 6779 14841 6791 14844
rect 6733 14835 6791 14841
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 7116 14844 7604 14872
rect 4706 14804 4712 14816
rect 3988 14776 4712 14804
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 7116 14804 7144 14844
rect 7466 14804 7472 14816
rect 5684 14776 7144 14804
rect 7427 14776 7472 14804
rect 5684 14764 5690 14776
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 7576 14804 7604 14844
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 10502 14872 10508 14884
rect 10192 14844 10508 14872
rect 10192 14832 10198 14844
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 22066 14872 22094 14912
rect 26142 14900 26148 14912
rect 26200 14900 26206 14952
rect 26694 14900 26700 14952
rect 26752 14940 26758 14952
rect 27157 14943 27215 14949
rect 27157 14940 27169 14943
rect 26752 14912 27169 14940
rect 26752 14900 26758 14912
rect 27157 14909 27169 14912
rect 27203 14909 27215 14943
rect 27157 14903 27215 14909
rect 27341 14943 27399 14949
rect 27341 14909 27353 14943
rect 27387 14909 27399 14943
rect 27341 14903 27399 14909
rect 13004 14844 22094 14872
rect 27356 14872 27384 14903
rect 28629 14875 28687 14881
rect 28629 14872 28641 14875
rect 27356 14844 28641 14872
rect 9766 14804 9772 14816
rect 7576 14776 9772 14804
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 10778 14804 10784 14816
rect 10100 14776 10784 14804
rect 10100 14764 10106 14776
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11238 14764 11244 14816
rect 11296 14804 11302 14816
rect 13004 14804 13032 14844
rect 28629 14841 28641 14844
rect 28675 14841 28687 14875
rect 28629 14835 28687 14841
rect 11296 14776 13032 14804
rect 11296 14764 11302 14776
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 15286 14804 15292 14816
rect 13872 14776 15292 14804
rect 13872 14764 13878 14776
rect 15286 14764 15292 14776
rect 15344 14804 15350 14816
rect 18414 14804 18420 14816
rect 15344 14776 18420 14804
rect 15344 14764 15350 14776
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 24762 14764 24768 14816
rect 24820 14804 24826 14816
rect 26329 14807 26387 14813
rect 26329 14804 26341 14807
rect 24820 14776 26341 14804
rect 24820 14764 24826 14776
rect 26329 14773 26341 14776
rect 26375 14773 26387 14807
rect 26329 14767 26387 14773
rect 26786 14764 26792 14816
rect 26844 14804 26850 14816
rect 27525 14807 27583 14813
rect 27525 14804 27537 14807
rect 26844 14776 27537 14804
rect 26844 14764 26850 14776
rect 27525 14773 27537 14776
rect 27571 14773 27583 14807
rect 27525 14767 27583 14773
rect 37829 14807 37887 14813
rect 37829 14773 37841 14807
rect 37875 14804 37887 14807
rect 37918 14804 37924 14816
rect 37875 14776 37924 14804
rect 37875 14773 37887 14776
rect 37829 14767 37887 14773
rect 37918 14764 37924 14776
rect 37976 14764 37982 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 4893 14603 4951 14609
rect 4893 14569 4905 14603
rect 4939 14600 4951 14603
rect 7190 14600 7196 14612
rect 4939 14572 7052 14600
rect 7151 14572 7196 14600
rect 4939 14569 4951 14572
rect 4893 14563 4951 14569
rect 4798 14532 4804 14544
rect 4172 14504 4804 14532
rect 1578 14464 1584 14476
rect 1539 14436 1584 14464
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 4172 14473 4200 14504
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 5442 14492 5448 14544
rect 5500 14492 5506 14544
rect 7024 14532 7052 14572
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 7834 14600 7840 14612
rect 7795 14572 7840 14600
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 8018 14560 8024 14612
rect 8076 14600 8082 14612
rect 9858 14600 9864 14612
rect 8076 14572 9864 14600
rect 8076 14560 8082 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 14645 14603 14703 14609
rect 10008 14572 14596 14600
rect 10008 14560 10014 14572
rect 8662 14532 8668 14544
rect 7024 14504 8668 14532
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 10410 14492 10416 14544
rect 10468 14532 10474 14544
rect 13357 14535 13415 14541
rect 10468 14504 11652 14532
rect 10468 14492 10474 14504
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14433 4215 14467
rect 4157 14427 4215 14433
rect 3344 14396 3372 14427
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 5460 14464 5488 14492
rect 5718 14464 5724 14476
rect 4304 14436 5488 14464
rect 5679 14436 5724 14464
rect 4304 14424 4310 14436
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 9125 14467 9183 14473
rect 6512 14436 9076 14464
rect 6512 14424 6518 14436
rect 4801 14399 4859 14405
rect 4801 14396 4813 14399
rect 3344 14368 4813 14396
rect 4801 14365 4813 14368
rect 4847 14396 4859 14399
rect 4890 14396 4896 14408
rect 4847 14368 4896 14396
rect 4847 14365 4859 14368
rect 4801 14359 4859 14365
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 5442 14396 5448 14408
rect 5403 14368 5448 14396
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 7616 14368 7757 14396
rect 7616 14356 7622 14368
rect 7745 14365 7757 14368
rect 7791 14396 7803 14399
rect 8018 14396 8024 14408
rect 7791 14368 8024 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14396 8447 14399
rect 8846 14396 8852 14408
rect 8435 14368 8852 14396
rect 8435 14365 8447 14368
rect 8389 14359 8447 14365
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14297 1915 14331
rect 3082 14300 5764 14328
rect 1857 14291 1915 14297
rect 1872 14260 1900 14291
rect 2590 14260 2596 14272
rect 1872 14232 2596 14260
rect 2590 14220 2596 14232
rect 2648 14260 2654 14272
rect 5626 14260 5632 14272
rect 2648 14232 5632 14260
rect 2648 14220 2654 14232
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 5736 14260 5764 14300
rect 6730 14288 6736 14340
rect 6788 14288 6794 14340
rect 8481 14331 8539 14337
rect 8481 14328 8493 14331
rect 7024 14300 8493 14328
rect 7024 14260 7052 14300
rect 8481 14297 8493 14300
rect 8527 14297 8539 14331
rect 8481 14291 8539 14297
rect 5736 14232 7052 14260
rect 7190 14220 7196 14272
rect 7248 14260 7254 14272
rect 8386 14260 8392 14272
rect 7248 14232 8392 14260
rect 7248 14220 7254 14232
rect 8386 14220 8392 14232
rect 8444 14260 8450 14272
rect 8588 14260 8616 14368
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 8444 14232 8616 14260
rect 9048 14260 9076 14436
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 11514 14464 11520 14476
rect 9171 14436 11520 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 11624 14464 11652 14504
rect 13357 14501 13369 14535
rect 13403 14532 13415 14535
rect 13906 14532 13912 14544
rect 13403 14504 13912 14532
rect 13403 14501 13415 14504
rect 13357 14495 13415 14501
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 14568 14532 14596 14572
rect 14645 14569 14657 14603
rect 14691 14600 14703 14603
rect 16758 14600 16764 14612
rect 14691 14572 16764 14600
rect 14691 14569 14703 14572
rect 14645 14563 14703 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 20622 14600 20628 14612
rect 18288 14572 19564 14600
rect 20583 14572 20628 14600
rect 18288 14560 18294 14572
rect 15102 14532 15108 14544
rect 14568 14504 15108 14532
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 15194 14464 15200 14476
rect 11624 14436 15200 14464
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15470 14464 15476 14476
rect 15431 14436 15476 14464
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15620 14436 15761 14464
rect 15620 14424 15626 14436
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 17405 14467 17463 14473
rect 17405 14433 17417 14467
rect 17451 14464 17463 14467
rect 18598 14464 18604 14476
rect 17451 14436 18604 14464
rect 17451 14433 17463 14436
rect 17405 14427 17463 14433
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 18966 14424 18972 14476
rect 19024 14464 19030 14476
rect 19429 14467 19487 14473
rect 19429 14464 19441 14467
rect 19024 14436 19441 14464
rect 19024 14424 19030 14436
rect 19429 14433 19441 14436
rect 19475 14433 19487 14467
rect 19429 14427 19487 14433
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 10836 14368 11161 14396
rect 10836 14356 10842 14368
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 9398 14328 9404 14340
rect 9359 14300 9404 14328
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 9490 14288 9496 14340
rect 9548 14328 9554 14340
rect 10704 14328 10732 14356
rect 11624 14328 11652 14359
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 14516 14368 14565 14396
rect 14516 14356 14522 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18693 14399 18751 14405
rect 18693 14396 18705 14399
rect 18196 14368 18705 14396
rect 18196 14356 18202 14368
rect 18693 14365 18705 14368
rect 18739 14365 18751 14399
rect 19536 14396 19564 14572
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 21266 14560 21272 14612
rect 21324 14600 21330 14612
rect 34514 14600 34520 14612
rect 21324 14572 34520 14600
rect 21324 14560 21330 14572
rect 34514 14560 34520 14572
rect 34572 14560 34578 14612
rect 35345 14603 35403 14609
rect 35345 14569 35357 14603
rect 35391 14600 35403 14603
rect 36538 14600 36544 14612
rect 35391 14572 36544 14600
rect 35391 14569 35403 14572
rect 35345 14563 35403 14569
rect 36538 14560 36544 14572
rect 36596 14560 36602 14612
rect 20073 14535 20131 14541
rect 20073 14501 20085 14535
rect 20119 14532 20131 14535
rect 20898 14532 20904 14544
rect 20119 14504 20904 14532
rect 20119 14501 20131 14504
rect 20073 14495 20131 14501
rect 20898 14492 20904 14504
rect 20956 14492 20962 14544
rect 21450 14492 21456 14544
rect 21508 14532 21514 14544
rect 21508 14504 24624 14532
rect 21508 14492 21514 14504
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14464 19671 14467
rect 20254 14464 20260 14476
rect 19659 14436 20260 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 22002 14464 22008 14476
rect 20456 14436 22008 14464
rect 20456 14396 20484 14436
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 24596 14473 24624 14504
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14433 24639 14467
rect 24762 14464 24768 14476
rect 24723 14436 24768 14464
rect 24581 14427 24639 14433
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 26694 14464 26700 14476
rect 26655 14436 26700 14464
rect 26694 14424 26700 14436
rect 26752 14424 26758 14476
rect 19536 14368 20484 14396
rect 20533 14399 20591 14405
rect 18693 14359 18751 14365
rect 20533 14365 20545 14399
rect 20579 14396 20591 14399
rect 21542 14396 21548 14408
rect 20579 14368 21548 14396
rect 20579 14365 20591 14368
rect 20533 14359 20591 14365
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 21729 14399 21787 14405
rect 21729 14365 21741 14399
rect 21775 14396 21787 14399
rect 21910 14396 21916 14408
rect 21775 14368 21916 14396
rect 21775 14365 21787 14368
rect 21729 14359 21787 14365
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 26142 14356 26148 14408
rect 26200 14396 26206 14408
rect 27525 14399 27583 14405
rect 27525 14396 27537 14399
rect 26200 14368 27537 14396
rect 26200 14356 26206 14368
rect 27525 14365 27537 14368
rect 27571 14365 27583 14399
rect 27982 14396 27988 14408
rect 27943 14368 27988 14396
rect 27525 14359 27583 14365
rect 27982 14356 27988 14368
rect 28040 14356 28046 14408
rect 34606 14356 34612 14408
rect 34664 14396 34670 14408
rect 35529 14399 35587 14405
rect 35529 14396 35541 14399
rect 34664 14368 35541 14396
rect 34664 14356 34670 14368
rect 35529 14365 35541 14368
rect 35575 14365 35587 14399
rect 35529 14359 35587 14365
rect 37274 14356 37280 14408
rect 37332 14396 37338 14408
rect 38013 14399 38071 14405
rect 38013 14396 38025 14399
rect 37332 14368 38025 14396
rect 37332 14356 37338 14368
rect 38013 14365 38025 14368
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 9548 14300 9890 14328
rect 10704 14300 11652 14328
rect 9548 14288 9554 14300
rect 11790 14288 11796 14340
rect 11848 14328 11854 14340
rect 11885 14331 11943 14337
rect 11885 14328 11897 14331
rect 11848 14300 11897 14328
rect 11848 14288 11854 14300
rect 11885 14297 11897 14300
rect 11931 14297 11943 14331
rect 11885 14291 11943 14297
rect 11974 14288 11980 14340
rect 12032 14328 12038 14340
rect 15565 14331 15623 14337
rect 12032 14300 12374 14328
rect 13648 14300 14596 14328
rect 12032 14288 12038 14300
rect 10318 14260 10324 14272
rect 9048 14232 10324 14260
rect 8444 14220 8450 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10410 14220 10416 14272
rect 10468 14260 10474 14272
rect 13648 14260 13676 14300
rect 10468 14232 13676 14260
rect 14568 14260 14596 14300
rect 15565 14297 15577 14331
rect 15611 14297 15623 14331
rect 15565 14291 15623 14297
rect 17497 14331 17555 14337
rect 17497 14297 17509 14331
rect 17543 14328 17555 14331
rect 17862 14328 17868 14340
rect 17543 14300 17868 14328
rect 17543 14297 17555 14300
rect 17497 14291 17555 14297
rect 15580 14260 15608 14291
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 18049 14331 18107 14337
rect 18049 14297 18061 14331
rect 18095 14328 18107 14331
rect 20346 14328 20352 14340
rect 18095 14300 20352 14328
rect 18095 14297 18107 14300
rect 18049 14291 18107 14297
rect 14568 14232 15608 14260
rect 10468 14220 10474 14232
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17770 14260 17776 14272
rect 17092 14232 17776 14260
rect 17092 14220 17098 14232
rect 17770 14220 17776 14232
rect 17828 14260 17834 14272
rect 18064 14260 18092 14291
rect 20346 14288 20352 14300
rect 20404 14288 20410 14340
rect 17828 14232 18092 14260
rect 17828 14220 17834 14232
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 18785 14263 18843 14269
rect 18785 14260 18797 14263
rect 18748 14232 18797 14260
rect 18748 14220 18754 14232
rect 18785 14229 18797 14232
rect 18831 14229 18843 14263
rect 18785 14223 18843 14229
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 21821 14263 21879 14269
rect 21821 14260 21833 14263
rect 20956 14232 21833 14260
rect 20956 14220 20962 14232
rect 21821 14229 21833 14232
rect 21867 14229 21879 14263
rect 21821 14223 21879 14229
rect 25225 14263 25283 14269
rect 25225 14229 25237 14263
rect 25271 14260 25283 14263
rect 26602 14260 26608 14272
rect 25271 14232 26608 14260
rect 25271 14229 25283 14232
rect 25225 14223 25283 14229
rect 26602 14220 26608 14232
rect 26660 14220 26666 14272
rect 27338 14260 27344 14272
rect 27299 14232 27344 14260
rect 27338 14220 27344 14232
rect 27396 14220 27402 14272
rect 28074 14260 28080 14272
rect 28035 14232 28080 14260
rect 28074 14220 28080 14232
rect 28132 14220 28138 14272
rect 38194 14260 38200 14272
rect 38155 14232 38200 14260
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 2774 14056 2780 14068
rect 1811 14028 2780 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 13446 14056 13452 14068
rect 4908 14028 13308 14056
rect 13407 14028 13452 14056
rect 2409 13991 2467 13997
rect 2409 13957 2421 13991
rect 2455 13988 2467 13991
rect 4908 13988 4936 14028
rect 6454 13988 6460 14000
rect 2455 13960 4936 13988
rect 5750 13960 6460 13988
rect 2455 13957 2467 13960
rect 2409 13951 2467 13957
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 6641 13991 6699 13997
rect 6641 13957 6653 13991
rect 6687 13988 6699 13991
rect 7374 13988 7380 14000
rect 6687 13960 7380 13988
rect 6687 13957 6699 13960
rect 6641 13951 6699 13957
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 7466 13948 7472 14000
rect 7524 13988 7530 14000
rect 9861 13991 9919 13997
rect 7524 13960 8602 13988
rect 7524 13948 7530 13960
rect 9861 13957 9873 13991
rect 9907 13988 9919 13991
rect 10042 13988 10048 14000
rect 9907 13960 10048 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 10042 13948 10048 13960
rect 10100 13948 10106 14000
rect 10410 13988 10416 14000
rect 10371 13960 10416 13988
rect 10410 13948 10416 13960
rect 10468 13948 10474 14000
rect 11054 13988 11060 14000
rect 11015 13960 11060 13988
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 12434 13948 12440 14000
rect 12492 13948 12498 14000
rect 13280 13988 13308 14028
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 15010 14056 15016 14068
rect 13740 14028 15016 14056
rect 13740 13988 13768 14028
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 15657 14059 15715 14065
rect 15657 14056 15669 14059
rect 15120 14028 15669 14056
rect 13280 13960 13768 13988
rect 14090 13948 14096 14000
rect 14148 13988 14154 14000
rect 14148 13960 14193 13988
rect 14148 13948 14154 13960
rect 14274 13948 14280 14000
rect 14332 13988 14338 14000
rect 15120 13988 15148 14028
rect 15657 14025 15669 14028
rect 15703 14025 15715 14059
rect 20530 14056 20536 14068
rect 15657 14019 15715 14025
rect 17144 14028 20536 14056
rect 14332 13960 15148 13988
rect 14332 13948 14338 13960
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 17034 13988 17040 14000
rect 15252 13960 15608 13988
rect 16995 13960 17040 13988
rect 15252 13948 15258 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 1581 13883 1639 13889
rect 1596 13852 1624 13883
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2823 13892 3065 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 3053 13889 3065 13892
rect 3099 13920 3111 13923
rect 4154 13920 4160 13932
rect 3099 13892 4160 13920
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 7190 13920 7196 13932
rect 7151 13892 7196 13920
rect 6549 13883 6607 13889
rect 2682 13852 2688 13864
rect 1596 13824 2688 13852
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 5258 13852 5264 13864
rect 4571 13824 5264 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 3234 13716 3240 13728
rect 3195 13688 3240 13716
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 4264 13716 4292 13815
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6270 13852 6276 13864
rect 6043 13824 6276 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 6564 13852 6592 13883
rect 7190 13880 7196 13892
rect 7248 13880 7254 13932
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 9548 13892 10333 13920
rect 9548 13880 9554 13892
rect 10321 13889 10333 13892
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10778 13920 10784 13932
rect 10560 13892 10784 13920
rect 10560 13880 10566 13892
rect 10778 13880 10784 13892
rect 10836 13920 10842 13932
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10836 13892 10977 13920
rect 10836 13880 10842 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 11698 13920 11704 13932
rect 11659 13892 11704 13920
rect 10965 13883 11023 13889
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 15580 13929 15608 13960
rect 17034 13948 17040 13960
rect 17092 13948 17098 14000
rect 17144 13997 17172 14028
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 22462 14056 22468 14068
rect 22204 14028 22468 14056
rect 17129 13991 17187 13997
rect 17129 13957 17141 13991
rect 17175 13957 17187 13991
rect 17129 13951 17187 13957
rect 17678 13948 17684 14000
rect 17736 13988 17742 14000
rect 18049 13991 18107 13997
rect 18049 13988 18061 13991
rect 17736 13960 18061 13988
rect 17736 13948 17742 13960
rect 18049 13957 18061 13960
rect 18095 13957 18107 13991
rect 18690 13988 18696 14000
rect 18651 13960 18696 13988
rect 18049 13951 18107 13957
rect 18690 13948 18696 13960
rect 18748 13948 18754 14000
rect 20349 13991 20407 13997
rect 20349 13957 20361 13991
rect 20395 13988 20407 13991
rect 22204 13988 22232 14028
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 26602 14056 26608 14068
rect 26563 14028 26608 14056
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 27157 14059 27215 14065
rect 27157 14025 27169 14059
rect 27203 14025 27215 14059
rect 27157 14019 27215 14025
rect 33689 14059 33747 14065
rect 33689 14025 33701 14059
rect 33735 14056 33747 14059
rect 34790 14056 34796 14068
rect 33735 14028 34796 14056
rect 33735 14025 33747 14028
rect 33689 14019 33747 14025
rect 26786 13988 26792 14000
rect 20395 13960 22232 13988
rect 25976 13960 26792 13988
rect 20395 13957 20407 13960
rect 20349 13951 20407 13957
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 20806 13920 20812 13932
rect 15565 13883 15623 13889
rect 17880 13892 18184 13920
rect 20767 13892 20812 13920
rect 7466 13852 7472 13864
rect 6564 13824 7472 13852
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 7834 13852 7840 13864
rect 7795 13824 7840 13852
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8113 13855 8171 13861
rect 8113 13821 8125 13855
rect 8159 13852 8171 13855
rect 8159 13824 9168 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 9140 13784 9168 13824
rect 9398 13812 9404 13864
rect 9456 13852 9462 13864
rect 10042 13852 10048 13864
rect 9456 13824 10048 13852
rect 9456 13812 9462 13824
rect 10042 13812 10048 13824
rect 10100 13812 10106 13864
rect 11974 13852 11980 13864
rect 11935 13824 11980 13852
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14642 13852 14648 13864
rect 14047 13824 14648 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15470 13852 15476 13864
rect 15059 13824 15476 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 17494 13812 17500 13864
rect 17552 13852 17558 13864
rect 17880 13852 17908 13892
rect 17552 13824 17908 13852
rect 18156 13852 18184 13892
rect 20806 13880 20812 13892
rect 20864 13880 20870 13932
rect 22370 13880 22376 13932
rect 22428 13920 22434 13932
rect 22925 13923 22983 13929
rect 22925 13920 22937 13923
rect 22428 13892 22937 13920
rect 22428 13880 22434 13892
rect 22925 13889 22937 13892
rect 22971 13889 22983 13923
rect 23566 13920 23572 13932
rect 23527 13892 23572 13920
rect 22925 13883 22983 13889
rect 23566 13880 23572 13892
rect 23624 13880 23630 13932
rect 25976 13929 26004 13960
rect 26786 13948 26792 13960
rect 26844 13948 26850 14000
rect 25961 13923 26019 13929
rect 25961 13889 25973 13923
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 26145 13923 26203 13929
rect 26145 13889 26157 13923
rect 26191 13920 26203 13923
rect 27172 13920 27200 14019
rect 34790 14016 34796 14028
rect 34848 14016 34854 14068
rect 27338 13920 27344 13932
rect 26191 13892 27200 13920
rect 27299 13892 27344 13920
rect 26191 13889 26203 13892
rect 26145 13883 26203 13889
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13889 27859 13923
rect 27801 13883 27859 13889
rect 27893 13923 27951 13929
rect 27893 13889 27905 13923
rect 27939 13920 27951 13923
rect 33873 13923 33931 13929
rect 33873 13920 33885 13923
rect 27939 13892 33885 13920
rect 27939 13889 27951 13892
rect 27893 13883 27951 13889
rect 33873 13889 33885 13892
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18156 13824 18613 13852
rect 17552 13812 17558 13824
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 18601 13815 18659 13821
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18840 13824 18889 13852
rect 18840 13812 18846 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 19702 13852 19708 13864
rect 19663 13824 19708 13852
rect 18877 13815 18935 13821
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 19889 13855 19947 13861
rect 19889 13821 19901 13855
rect 19935 13852 19947 13855
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 19935 13824 20913 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 22152 13824 22293 13852
rect 22152 13812 22158 13824
rect 22281 13821 22293 13824
rect 22327 13821 22339 13855
rect 22462 13852 22468 13864
rect 22423 13824 22468 13852
rect 22281 13815 22339 13821
rect 22462 13812 22468 13824
rect 22520 13812 22526 13864
rect 26602 13812 26608 13864
rect 26660 13852 26666 13864
rect 27816 13852 27844 13883
rect 26660 13824 27844 13852
rect 26660 13812 26666 13824
rect 10226 13784 10232 13796
rect 6788 13756 7420 13784
rect 9140 13756 10232 13784
rect 6788 13744 6794 13756
rect 4614 13716 4620 13728
rect 4264 13688 4620 13716
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7285 13719 7343 13725
rect 7285 13716 7297 13719
rect 7248 13688 7297 13716
rect 7248 13676 7254 13688
rect 7285 13685 7297 13688
rect 7331 13685 7343 13719
rect 7392 13716 7420 13756
rect 10226 13744 10232 13756
rect 10284 13744 10290 13796
rect 17218 13784 17224 13796
rect 13372 13756 17224 13784
rect 13372 13716 13400 13756
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 20990 13784 20996 13796
rect 19306 13756 20996 13784
rect 7392 13688 13400 13716
rect 7285 13679 7343 13685
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 15102 13716 15108 13728
rect 13964 13688 15108 13716
rect 13964 13676 13970 13688
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 16114 13676 16120 13728
rect 16172 13716 16178 13728
rect 19306 13716 19334 13756
rect 20990 13744 20996 13756
rect 21048 13744 21054 13796
rect 21082 13744 21088 13796
rect 21140 13784 21146 13796
rect 23290 13784 23296 13796
rect 21140 13756 23296 13784
rect 21140 13744 21146 13756
rect 23290 13744 23296 13756
rect 23348 13744 23354 13796
rect 16172 13688 19334 13716
rect 16172 13676 16178 13688
rect 19702 13676 19708 13728
rect 19760 13716 19766 13728
rect 22922 13716 22928 13728
rect 19760 13688 22928 13716
rect 19760 13676 19766 13688
rect 22922 13676 22928 13688
rect 22980 13676 22986 13728
rect 23382 13716 23388 13728
rect 23343 13688 23388 13716
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 1844 13515 1902 13521
rect 1844 13481 1856 13515
rect 1890 13512 1902 13515
rect 2958 13512 2964 13524
rect 1890 13484 2964 13512
rect 1890 13481 1902 13484
rect 1844 13475 1902 13481
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 3326 13512 3332 13524
rect 3239 13484 3332 13512
rect 3326 13472 3332 13484
rect 3384 13512 3390 13524
rect 5350 13512 5356 13524
rect 3384 13484 5356 13512
rect 3384 13472 3390 13484
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 9490 13512 9496 13524
rect 6144 13484 9496 13512
rect 6144 13472 6150 13484
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10008 13484 10885 13512
rect 10008 13472 10014 13484
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 10873 13475 10931 13481
rect 11974 13472 11980 13524
rect 12032 13512 12038 13524
rect 14458 13512 14464 13524
rect 12032 13484 14464 13512
rect 12032 13472 12038 13484
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 18230 13512 18236 13524
rect 14568 13484 18236 13512
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 9030 13444 9036 13456
rect 7607 13416 9036 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 13630 13404 13636 13456
rect 13688 13444 13694 13456
rect 14568 13444 14596 13484
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19889 13515 19947 13521
rect 19889 13481 19901 13515
rect 19935 13512 19947 13515
rect 20070 13512 20076 13524
rect 19935 13484 20076 13512
rect 19935 13481 19947 13484
rect 19889 13475 19947 13481
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20530 13472 20536 13524
rect 20588 13512 20594 13524
rect 21637 13515 21695 13521
rect 21637 13512 21649 13515
rect 20588 13484 21649 13512
rect 20588 13472 20594 13484
rect 21637 13481 21649 13484
rect 21683 13481 21695 13515
rect 22462 13512 22468 13524
rect 22423 13484 22468 13512
rect 21637 13475 21695 13481
rect 22462 13472 22468 13484
rect 22520 13472 22526 13524
rect 26786 13512 26792 13524
rect 26747 13484 26792 13512
rect 26786 13472 26792 13484
rect 26844 13472 26850 13524
rect 13688 13416 14596 13444
rect 13688 13404 13694 13416
rect 18046 13404 18052 13456
rect 18104 13444 18110 13456
rect 20438 13444 20444 13456
rect 18104 13416 20444 13444
rect 18104 13404 18110 13416
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 26234 13444 26240 13456
rect 20548 13416 26240 13444
rect 1578 13376 1584 13388
rect 1491 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13376 1642 13388
rect 4614 13376 4620 13388
rect 1636 13348 4620 13376
rect 1636 13336 1642 13348
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 8938 13376 8944 13388
rect 6604 13348 8944 13376
rect 6604 13336 6610 13348
rect 8938 13336 8944 13348
rect 8996 13336 9002 13388
rect 9122 13376 9128 13388
rect 9083 13348 9128 13376
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 11238 13376 11244 13388
rect 9456 13348 11244 13376
rect 9456 13336 9462 13348
rect 11238 13336 11244 13348
rect 11296 13336 11302 13388
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11698 13376 11704 13388
rect 11379 13348 11704 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 14366 13376 14372 13388
rect 12676 13348 13124 13376
rect 14327 13348 14372 13376
rect 12676 13336 12682 13348
rect 13096 13320 13124 13348
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 15378 13376 15384 13388
rect 15339 13348 15384 13376
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 16577 13379 16635 13385
rect 16577 13345 16589 13379
rect 16623 13376 16635 13379
rect 16666 13376 16672 13388
rect 16623 13348 16672 13376
rect 16623 13345 16635 13348
rect 16577 13339 16635 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16942 13376 16948 13388
rect 16903 13348 16948 13376
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 20548 13376 20576 13416
rect 26234 13404 26240 13416
rect 26292 13444 26298 13456
rect 27246 13444 27252 13456
rect 26292 13416 27252 13444
rect 26292 13404 26298 13416
rect 27246 13404 27252 13416
rect 27304 13404 27310 13456
rect 17092 13348 20576 13376
rect 20625 13379 20683 13385
rect 17092 13336 17098 13348
rect 20625 13345 20637 13379
rect 20671 13376 20683 13379
rect 20898 13376 20904 13388
rect 20671 13348 20904 13376
rect 20671 13345 20683 13348
rect 20625 13339 20683 13345
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 21085 13379 21143 13385
rect 21085 13345 21097 13379
rect 21131 13376 21143 13379
rect 22830 13376 22836 13388
rect 21131 13348 22836 13376
rect 21131 13345 21143 13348
rect 21085 13339 21143 13345
rect 22830 13336 22836 13348
rect 22888 13336 22894 13388
rect 28074 13376 28080 13388
rect 26344 13348 28080 13376
rect 3970 13308 3976 13320
rect 3931 13280 3976 13308
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 5442 13308 5448 13320
rect 4212 13280 5448 13308
rect 4212 13268 4218 13280
rect 5442 13268 5448 13280
rect 5500 13308 5506 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5500 13280 5825 13308
rect 5500 13268 5506 13280
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 3082 13212 4016 13240
rect 3988 13184 4016 13212
rect 4614 13200 4620 13252
rect 4672 13240 4678 13252
rect 4709 13243 4767 13249
rect 4709 13240 4721 13243
rect 4672 13212 4721 13240
rect 4672 13200 4678 13212
rect 4709 13209 4721 13212
rect 4755 13209 4767 13243
rect 4709 13203 4767 13209
rect 3970 13132 3976 13184
rect 4028 13132 4034 13184
rect 5828 13172 5856 13271
rect 7190 13268 7196 13320
rect 7248 13268 7254 13320
rect 8386 13308 8392 13320
rect 8347 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13268 8450 13320
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 13136 13280 13369 13308
rect 13136 13268 13142 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13446 13268 13452 13320
rect 13504 13308 13510 13320
rect 15841 13311 15899 13317
rect 13504 13280 13952 13308
rect 13504 13268 13510 13280
rect 5994 13200 6000 13252
rect 6052 13240 6058 13252
rect 6089 13243 6147 13249
rect 6089 13240 6101 13243
rect 6052 13212 6101 13240
rect 6052 13200 6058 13212
rect 6089 13209 6101 13212
rect 6135 13209 6147 13243
rect 6089 13203 6147 13209
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 8260 13212 8708 13240
rect 8260 13200 8266 13212
rect 7098 13172 7104 13184
rect 5828 13144 7104 13172
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 8680 13172 8708 13212
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9088 13212 9413 13240
rect 9088 13200 9094 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 9508 13212 9890 13240
rect 9508 13172 9536 13212
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 11609 13243 11667 13249
rect 11609 13240 11621 13243
rect 11572 13212 11621 13240
rect 11572 13200 11578 13212
rect 11609 13209 11621 13212
rect 11655 13209 11667 13243
rect 11609 13203 11667 13209
rect 12066 13200 12072 13252
rect 12124 13200 12130 13252
rect 13538 13200 13544 13252
rect 13596 13240 13602 13252
rect 13924 13240 13952 13280
rect 15841 13277 15853 13311
rect 15887 13308 15899 13311
rect 16114 13308 16120 13320
rect 15887 13280 16120 13308
rect 15887 13277 15899 13280
rect 15841 13271 15899 13277
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 18598 13308 18604 13320
rect 18559 13280 18604 13308
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 19702 13308 19708 13320
rect 18840 13280 19708 13308
rect 18840 13268 18846 13280
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 14461 13243 14519 13249
rect 14461 13240 14473 13243
rect 13596 13212 13860 13240
rect 13924 13212 14473 13240
rect 13596 13200 13602 13212
rect 8680 13144 9536 13172
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 11238 13172 11244 13184
rect 9640 13144 11244 13172
rect 9640 13132 9646 13144
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 13722 13172 13728 13184
rect 12400 13144 13728 13172
rect 12400 13132 12406 13144
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 13832 13172 13860 13212
rect 14461 13209 14473 13212
rect 14507 13209 14519 13243
rect 16669 13243 16727 13249
rect 14461 13203 14519 13209
rect 14660 13212 16068 13240
rect 14660 13172 14688 13212
rect 13832 13144 14688 13172
rect 15102 13132 15108 13184
rect 15160 13172 15166 13184
rect 15933 13175 15991 13181
rect 15933 13172 15945 13175
rect 15160 13144 15945 13172
rect 15160 13132 15166 13144
rect 15933 13141 15945 13144
rect 15979 13141 15991 13175
rect 16040 13172 16068 13212
rect 16669 13209 16681 13243
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 17865 13243 17923 13249
rect 17865 13209 17877 13243
rect 17911 13240 17923 13243
rect 19812 13240 19840 13271
rect 20162 13268 20168 13320
rect 20220 13308 20226 13320
rect 20441 13311 20499 13317
rect 20441 13308 20453 13311
rect 20220 13280 20453 13308
rect 20220 13268 20226 13280
rect 20441 13277 20453 13280
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 20864 13280 21557 13308
rect 20864 13268 20870 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13308 22707 13311
rect 23382 13308 23388 13320
rect 22695 13280 23388 13308
rect 22695 13277 22707 13280
rect 22649 13271 22707 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23934 13308 23940 13320
rect 23895 13280 23940 13308
rect 23934 13268 23940 13280
rect 23992 13268 23998 13320
rect 25866 13268 25872 13320
rect 25924 13308 25930 13320
rect 26344 13317 26372 13348
rect 28074 13336 28080 13348
rect 28132 13336 28138 13388
rect 26145 13311 26203 13317
rect 26145 13308 26157 13311
rect 25924 13280 26157 13308
rect 25924 13268 25930 13280
rect 26145 13277 26157 13280
rect 26191 13277 26203 13311
rect 26145 13271 26203 13277
rect 26329 13311 26387 13317
rect 26329 13277 26341 13311
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 27246 13268 27252 13320
rect 27304 13308 27310 13320
rect 27304 13280 27349 13308
rect 27304 13268 27310 13280
rect 34790 13268 34796 13320
rect 34848 13308 34854 13320
rect 38013 13311 38071 13317
rect 38013 13308 38025 13311
rect 34848 13280 38025 13308
rect 34848 13268 34854 13280
rect 38013 13277 38025 13280
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 20254 13240 20260 13252
rect 17911 13212 19334 13240
rect 19812 13212 20260 13240
rect 17911 13209 17923 13212
rect 17865 13203 17923 13209
rect 16684 13172 16712 13203
rect 17954 13172 17960 13184
rect 16040 13144 16712 13172
rect 17915 13144 17960 13172
rect 15933 13135 15991 13141
rect 17954 13132 17960 13144
rect 18012 13132 18018 13184
rect 18690 13172 18696 13184
rect 18651 13144 18696 13172
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 19306 13172 19334 13212
rect 20254 13200 20260 13212
rect 20312 13200 20318 13252
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 22738 13240 22744 13252
rect 20404 13212 22744 13240
rect 20404 13200 20410 13212
rect 22738 13200 22744 13212
rect 22796 13200 22802 13252
rect 37274 13240 37280 13252
rect 23768 13212 37280 13240
rect 20714 13172 20720 13184
rect 19306 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 20990 13132 20996 13184
rect 21048 13172 21054 13184
rect 23658 13172 23664 13184
rect 21048 13144 23664 13172
rect 21048 13132 21054 13144
rect 23658 13132 23664 13144
rect 23716 13132 23722 13184
rect 23768 13181 23796 13212
rect 37274 13200 37280 13212
rect 37332 13200 37338 13252
rect 23753 13175 23811 13181
rect 23753 13141 23765 13175
rect 23799 13141 23811 13175
rect 27338 13172 27344 13184
rect 27299 13144 27344 13172
rect 23753 13135 23811 13141
rect 27338 13132 27344 13144
rect 27396 13132 27402 13184
rect 38194 13172 38200 13184
rect 38155 13144 38200 13172
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 3326 12968 3332 12980
rect 1872 12940 3332 12968
rect 1872 12909 1900 12940
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 4172 12940 6009 12968
rect 1857 12903 1915 12909
rect 1857 12869 1869 12903
rect 1903 12869 1915 12903
rect 4062 12900 4068 12912
rect 3082 12872 4068 12900
rect 1857 12863 1915 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 4172 12832 4200 12940
rect 5997 12937 6009 12940
rect 6043 12968 6055 12971
rect 6086 12968 6092 12980
rect 6043 12940 6092 12968
rect 6043 12937 6055 12940
rect 5997 12931 6055 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 6687 12940 9536 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 6822 12900 6828 12912
rect 5750 12872 6828 12900
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 7926 12860 7932 12912
rect 7984 12860 7990 12912
rect 9214 12900 9220 12912
rect 9175 12872 9220 12900
rect 9214 12860 9220 12872
rect 9272 12860 9278 12912
rect 3252 12804 4200 12832
rect 1578 12764 1584 12776
rect 1539 12736 1584 12764
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 3252 12628 3280 12804
rect 5994 12792 6000 12844
rect 6052 12832 6058 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6052 12804 6561 12832
rect 6052 12792 6058 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 7156 12804 7205 12832
rect 7156 12792 7162 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9508 12832 9536 12940
rect 10060 12940 14228 12968
rect 10060 12912 10088 12940
rect 14200 12912 14228 12940
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 15102 12968 15108 12980
rect 14792 12940 15108 12968
rect 14792 12928 14798 12940
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17184 12940 19840 12968
rect 17184 12928 17190 12940
rect 9674 12900 9680 12912
rect 9635 12872 9680 12900
rect 9674 12860 9680 12872
rect 9732 12900 9738 12912
rect 10042 12900 10048 12912
rect 9732 12872 10048 12900
rect 9732 12860 9738 12872
rect 10042 12860 10048 12872
rect 10100 12860 10106 12912
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 13722 12900 13728 12912
rect 11296 12872 12466 12900
rect 13683 12872 13728 12900
rect 11296 12860 11302 12872
rect 13722 12860 13728 12872
rect 13780 12860 13786 12912
rect 14182 12900 14188 12912
rect 14095 12872 14188 12900
rect 14182 12860 14188 12872
rect 14240 12860 14246 12912
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12900 15807 12903
rect 18690 12900 18696 12912
rect 15795 12872 18460 12900
rect 18651 12872 18696 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 11698 12832 11704 12844
rect 9180 12804 9444 12832
rect 9508 12804 11560 12832
rect 11659 12804 11704 12832
rect 9180 12792 9186 12804
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 3384 12736 3429 12764
rect 3384 12724 3390 12736
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4249 12767 4307 12773
rect 4249 12764 4261 12767
rect 4212 12736 4261 12764
rect 4212 12724 4218 12736
rect 4249 12733 4261 12736
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5534 12764 5540 12776
rect 4571 12736 5540 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12764 7527 12767
rect 8662 12764 8668 12776
rect 7515 12736 8668 12764
rect 7515 12733 7527 12736
rect 7469 12727 7527 12733
rect 8662 12724 8668 12736
rect 8720 12764 8726 12776
rect 9306 12764 9312 12776
rect 8720 12736 9312 12764
rect 8720 12724 8726 12736
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 9416 12764 9444 12804
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 9416 12736 10517 12764
rect 10505 12733 10517 12736
rect 10551 12764 10563 12767
rect 11238 12764 11244 12776
rect 10551 12736 11244 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 8938 12656 8944 12708
rect 8996 12696 9002 12708
rect 9950 12696 9956 12708
rect 8996 12668 9956 12696
rect 8996 12656 9002 12668
rect 9950 12656 9956 12668
rect 10008 12656 10014 12708
rect 2096 12600 3280 12628
rect 2096 12588 2102 12600
rect 4982 12588 4988 12640
rect 5040 12628 5046 12640
rect 7282 12628 7288 12640
rect 5040 12600 7288 12628
rect 5040 12588 5046 12600
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 9122 12628 9128 12640
rect 7892 12600 9128 12628
rect 7892 12588 7898 12600
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 11146 12628 11152 12640
rect 9548 12600 11152 12628
rect 9548 12588 9554 12600
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11532 12628 11560 12804
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 17218 12832 17224 12844
rect 17179 12804 17224 12832
rect 17218 12792 17224 12804
rect 17276 12832 17282 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17276 12804 17877 12832
rect 17276 12792 17282 12804
rect 17865 12801 17877 12804
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12764 12035 12767
rect 12618 12764 12624 12776
rect 12023 12736 12624 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12618 12724 12624 12736
rect 12676 12724 12682 12776
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14056 12736 14933 12764
rect 14056 12724 14062 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 15654 12764 15660 12776
rect 15615 12736 15660 12764
rect 14921 12727 14979 12733
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 17678 12764 17684 12776
rect 16132 12736 17684 12764
rect 14090 12696 14096 12708
rect 13004 12668 14096 12696
rect 13004 12628 13032 12668
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 11532 12600 13032 12628
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 16132 12628 16160 12736
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 16209 12699 16267 12705
rect 16209 12665 16221 12699
rect 16255 12696 16267 12699
rect 17218 12696 17224 12708
rect 16255 12668 17224 12696
rect 16255 12665 16267 12668
rect 16209 12659 16267 12665
rect 17218 12656 17224 12668
rect 17276 12656 17282 12708
rect 17696 12696 17724 12724
rect 18432 12696 18460 12872
rect 18690 12860 18696 12872
rect 18748 12860 18754 12912
rect 19812 12832 19840 12940
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 23934 12968 23940 12980
rect 20036 12940 23940 12968
rect 20036 12928 20042 12940
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 22738 12900 22744 12912
rect 22699 12872 22744 12900
rect 22738 12860 22744 12872
rect 22796 12860 22802 12912
rect 23382 12900 23388 12912
rect 23343 12872 23388 12900
rect 23382 12860 23388 12872
rect 23440 12860 23446 12912
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 19444 12804 19748 12832
rect 19812 12804 20085 12832
rect 18601 12767 18659 12773
rect 18601 12733 18613 12767
rect 18647 12764 18659 12767
rect 18782 12764 18788 12776
rect 18647 12736 18788 12764
rect 18647 12733 18659 12736
rect 18601 12727 18659 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 18966 12724 18972 12776
rect 19024 12764 19030 12776
rect 19444 12764 19472 12804
rect 19610 12764 19616 12776
rect 19024 12736 19472 12764
rect 19571 12736 19616 12764
rect 19024 12724 19030 12736
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19720 12764 19748 12804
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20714 12832 20720 12844
rect 20627 12804 20720 12832
rect 20073 12795 20131 12801
rect 20714 12792 20720 12804
rect 20772 12832 20778 12844
rect 21818 12832 21824 12844
rect 20772 12804 21824 12832
rect 20772 12792 20778 12804
rect 21818 12792 21824 12804
rect 21876 12792 21882 12844
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12801 22063 12835
rect 22649 12835 22707 12841
rect 22649 12832 22661 12835
rect 22005 12795 22063 12801
rect 22112 12804 22661 12832
rect 22020 12764 22048 12795
rect 19720 12736 22048 12764
rect 20346 12696 20352 12708
rect 17696 12668 18368 12696
rect 18432 12668 20352 12696
rect 17310 12628 17316 12640
rect 15068 12600 16160 12628
rect 17271 12600 17316 12628
rect 15068 12588 15074 12600
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 17954 12628 17960 12640
rect 17915 12600 17960 12628
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18340 12628 18368 12668
rect 20346 12656 20352 12668
rect 20404 12656 20410 12708
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 22112 12696 22140 12804
rect 22649 12801 22661 12804
rect 22695 12801 22707 12835
rect 23290 12832 23296 12844
rect 23251 12804 23296 12832
rect 22649 12795 22707 12801
rect 23290 12792 23296 12804
rect 23348 12792 23354 12844
rect 38286 12832 38292 12844
rect 38247 12804 38292 12832
rect 38286 12792 38292 12804
rect 38344 12792 38350 12844
rect 20496 12668 22140 12696
rect 20496 12656 20502 12668
rect 19978 12628 19984 12640
rect 18340 12600 19984 12628
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20165 12631 20223 12637
rect 20165 12597 20177 12631
rect 20211 12628 20223 12631
rect 20622 12628 20628 12640
rect 20211 12600 20628 12628
rect 20211 12597 20223 12600
rect 20165 12591 20223 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 20809 12631 20867 12637
rect 20809 12597 20821 12631
rect 20855 12628 20867 12631
rect 20990 12628 20996 12640
rect 20855 12600 20996 12628
rect 20855 12597 20867 12600
rect 20809 12591 20867 12597
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22152 12600 22197 12628
rect 22152 12588 22158 12600
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 22830 12628 22836 12640
rect 22612 12600 22836 12628
rect 22612 12588 22618 12600
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 38102 12628 38108 12640
rect 38063 12600 38108 12628
rect 38102 12588 38108 12600
rect 38160 12588 38166 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 3142 12384 3148 12436
rect 3200 12424 3206 12436
rect 3326 12424 3332 12436
rect 3200 12396 3332 12424
rect 3200 12384 3206 12396
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 4062 12424 4068 12436
rect 3896 12396 4068 12424
rect 1578 12248 1584 12300
rect 1636 12288 1642 12300
rect 1673 12291 1731 12297
rect 1673 12288 1685 12291
rect 1636 12260 1685 12288
rect 1636 12248 1642 12260
rect 1673 12257 1685 12260
rect 1719 12257 1731 12291
rect 1673 12251 1731 12257
rect 3896 12220 3924 12396
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 5442 12424 5448 12436
rect 4764 12396 5448 12424
rect 4764 12384 4770 12396
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 8481 12427 8539 12433
rect 8481 12424 8493 12427
rect 5920 12396 8493 12424
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 5920 12288 5948 12396
rect 8481 12393 8493 12396
rect 8527 12393 8539 12427
rect 8481 12387 8539 12393
rect 8496 12356 8524 12387
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 10686 12424 10692 12436
rect 9364 12396 10692 12424
rect 9364 12384 9370 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 12710 12384 12716 12436
rect 12768 12424 12774 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 12768 12396 13001 12424
rect 12768 12384 12774 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 13538 12424 13544 12436
rect 13499 12396 13544 12424
rect 12989 12387 13047 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 13780 12396 17909 12424
rect 13780 12384 13786 12396
rect 16022 12356 16028 12368
rect 8496 12328 11376 12356
rect 15983 12328 16028 12356
rect 7006 12288 7012 12300
rect 4304 12260 5948 12288
rect 6967 12260 7012 12288
rect 4304 12248 4310 12260
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 8018 12288 8024 12300
rect 7156 12260 8024 12288
rect 7156 12248 7162 12260
rect 8018 12248 8024 12260
rect 8076 12288 8082 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 8076 12260 9873 12288
rect 8076 12248 8082 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 11238 12288 11244 12300
rect 11199 12260 11244 12288
rect 9861 12251 9919 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11348 12288 11376 12328
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 16574 12316 16580 12368
rect 16632 12356 16638 12368
rect 16632 12328 17816 12356
rect 16632 12316 16638 12328
rect 14090 12288 14096 12300
rect 11348 12260 14096 12288
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 16040 12288 16068 12316
rect 14608 12260 16068 12288
rect 14608 12248 14614 12260
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 16908 12260 17693 12288
rect 16908 12248 16914 12260
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3896 12192 3985 12220
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 5350 12180 5356 12232
rect 5408 12180 5414 12232
rect 6730 12220 6736 12232
rect 6691 12192 6736 12220
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 8628 12192 10180 12220
rect 8628 12180 8634 12192
rect 1949 12155 2007 12161
rect 1949 12121 1961 12155
rect 1995 12121 2007 12155
rect 4154 12152 4160 12164
rect 3174 12124 4160 12152
rect 1949 12115 2007 12121
rect 1964 12084 1992 12115
rect 4154 12112 4160 12124
rect 4212 12112 4218 12164
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 4304 12124 4349 12152
rect 4304 12112 4310 12124
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 9030 12152 9036 12164
rect 5592 12124 6960 12152
rect 8234 12124 9036 12152
rect 5592 12112 5598 12124
rect 3234 12084 3240 12096
rect 1964 12056 3240 12084
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 3418 12084 3424 12096
rect 3379 12056 3424 12084
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 3568 12056 5733 12084
rect 3568 12044 3574 12056
rect 5721 12053 5733 12056
rect 5767 12053 5779 12087
rect 6932 12084 6960 12124
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 9125 12155 9183 12161
rect 9125 12121 9137 12155
rect 9171 12152 9183 12155
rect 9766 12152 9772 12164
rect 9171 12124 9772 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9766 12112 9772 12124
rect 9824 12152 9830 12164
rect 10042 12152 10048 12164
rect 9824 12124 10048 12152
rect 9824 12112 9830 12124
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 10152 12152 10180 12192
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 10284 12192 10609 12220
rect 10284 12180 10290 12192
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 13412 12192 13737 12220
rect 13412 12180 13418 12192
rect 13725 12189 13737 12192
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 14056 12192 14289 12220
rect 14056 12180 14062 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 16390 12220 16396 12232
rect 14277 12183 14335 12189
rect 15948 12192 16396 12220
rect 11238 12152 11244 12164
rect 10152 12124 11244 12152
rect 11238 12112 11244 12124
rect 11296 12112 11302 12164
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 11517 12155 11575 12161
rect 11517 12152 11529 12155
rect 11480 12124 11529 12152
rect 11480 12112 11486 12124
rect 11517 12121 11529 12124
rect 11563 12121 11575 12155
rect 11517 12115 11575 12121
rect 11790 12112 11796 12164
rect 11848 12152 11854 12164
rect 11848 12124 11928 12152
rect 11848 12112 11854 12124
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 6932 12056 10701 12084
rect 5721 12047 5779 12053
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 11900 12084 11928 12124
rect 12250 12112 12256 12164
rect 12308 12112 12314 12164
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 12952 12124 14565 12152
rect 12952 12112 12958 12124
rect 14553 12121 14565 12124
rect 14599 12121 14611 12155
rect 14553 12115 14611 12121
rect 13906 12084 13912 12096
rect 11900 12056 13912 12084
rect 10689 12047 10747 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14568 12084 14596 12115
rect 15010 12112 15016 12164
rect 15068 12112 15074 12164
rect 15948 12084 15976 12192
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 17788 12220 17816 12328
rect 17881 12297 17909 12396
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 18196 12396 21220 12424
rect 18196 12384 18202 12396
rect 19889 12359 19947 12365
rect 19889 12325 19901 12359
rect 19935 12356 19947 12359
rect 20530 12356 20536 12368
rect 19935 12328 20536 12356
rect 19935 12325 19947 12328
rect 19889 12319 19947 12325
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 21192 12356 21220 12396
rect 21266 12384 21272 12436
rect 21324 12424 21330 12436
rect 22649 12427 22707 12433
rect 22649 12424 22661 12427
rect 21324 12396 22661 12424
rect 21324 12384 21330 12396
rect 22649 12393 22661 12396
rect 22695 12393 22707 12427
rect 23290 12424 23296 12436
rect 23251 12396 23296 12424
rect 22649 12387 22707 12393
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 21192 12328 23888 12356
rect 17865 12291 17923 12297
rect 17865 12257 17877 12291
rect 17911 12257 17923 12291
rect 17865 12251 17923 12257
rect 20898 12248 20904 12300
rect 20956 12288 20962 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 20956 12260 22017 12288
rect 20956 12248 20962 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 17788 12192 18337 12220
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 21910 12220 21916 12232
rect 21871 12192 21916 12220
rect 18325 12183 18383 12189
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 22554 12220 22560 12232
rect 22515 12192 22560 12220
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 23198 12220 23204 12232
rect 23159 12192 23204 12220
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 23860 12229 23888 12328
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 29733 12223 29791 12229
rect 29733 12189 29745 12223
rect 29779 12220 29791 12223
rect 38102 12220 38108 12232
rect 29779 12192 38108 12220
rect 29779 12189 29791 12192
rect 29733 12183 29791 12189
rect 38102 12180 38108 12192
rect 38160 12180 38166 12232
rect 16206 12112 16212 12164
rect 16264 12152 16270 12164
rect 16577 12155 16635 12161
rect 16577 12152 16589 12155
rect 16264 12124 16589 12152
rect 16264 12112 16270 12124
rect 16500 12096 16528 12124
rect 16577 12121 16589 12124
rect 16623 12121 16635 12155
rect 16577 12115 16635 12121
rect 16666 12112 16672 12164
rect 16724 12152 16730 12164
rect 17218 12152 17224 12164
rect 16724 12124 16769 12152
rect 17179 12124 17224 12152
rect 16724 12112 16730 12124
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 19705 12155 19763 12161
rect 19705 12121 19717 12155
rect 19751 12152 19763 12155
rect 19978 12152 19984 12164
rect 19751 12124 19984 12152
rect 19751 12121 19763 12124
rect 19705 12115 19763 12121
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 20438 12152 20444 12164
rect 20399 12124 20444 12152
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 20533 12155 20591 12161
rect 20533 12121 20545 12155
rect 20579 12152 20591 12155
rect 21266 12152 21272 12164
rect 20579 12124 21272 12152
rect 20579 12121 20591 12124
rect 20533 12115 20591 12121
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 21453 12155 21511 12161
rect 21453 12121 21465 12155
rect 21499 12121 21511 12155
rect 21453 12115 21511 12121
rect 14568 12056 15976 12084
rect 16482 12044 16488 12096
rect 16540 12044 16546 12096
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 20806 12084 20812 12096
rect 16816 12056 20812 12084
rect 16816 12044 16822 12056
rect 20806 12044 20812 12056
rect 20864 12044 20870 12096
rect 21082 12044 21088 12096
rect 21140 12084 21146 12096
rect 21468 12084 21496 12115
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 29825 12155 29883 12161
rect 29825 12152 29837 12155
rect 21600 12124 29837 12152
rect 21600 12112 21606 12124
rect 29825 12121 29837 12124
rect 29871 12121 29883 12155
rect 29825 12115 29883 12121
rect 21726 12084 21732 12096
rect 21140 12056 21732 12084
rect 21140 12044 21146 12056
rect 21726 12044 21732 12056
rect 21784 12044 21790 12096
rect 22462 12044 22468 12096
rect 22520 12084 22526 12096
rect 23937 12087 23995 12093
rect 23937 12084 23949 12087
rect 22520 12056 23949 12084
rect 22520 12044 22526 12056
rect 23937 12053 23949 12056
rect 23983 12053 23995 12087
rect 23937 12047 23995 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 1946 11840 1952 11892
rect 2004 11880 2010 11892
rect 3602 11880 3608 11892
rect 2004 11852 3608 11880
rect 2004 11840 2010 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4212 11852 5856 11880
rect 4212 11840 4218 11852
rect 1854 11812 1860 11824
rect 1815 11784 1860 11812
rect 1854 11772 1860 11784
rect 1912 11772 1918 11824
rect 4614 11812 4620 11824
rect 4264 11784 4620 11812
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 4264 11753 4292 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 4249 11747 4307 11753
rect 2990 11716 4200 11744
rect 1210 11636 1216 11688
rect 1268 11676 1274 11688
rect 1946 11676 1952 11688
rect 1268 11648 1952 11676
rect 1268 11636 1274 11648
rect 1946 11636 1952 11648
rect 2004 11676 2010 11688
rect 3510 11676 3516 11688
rect 2004 11648 3516 11676
rect 2004 11636 2010 11648
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3660 11648 3705 11676
rect 3660 11636 3666 11648
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 3510 11540 3516 11552
rect 2372 11512 3516 11540
rect 2372 11500 2378 11512
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 4172 11540 4200 11716
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 4522 11676 4528 11688
rect 4483 11648 4528 11676
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 5644 11608 5672 11730
rect 5828 11676 5856 11852
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9088 11852 9904 11880
rect 9088 11840 9094 11852
rect 6730 11772 6736 11824
rect 6788 11812 6794 11824
rect 7834 11812 7840 11824
rect 6788 11784 7840 11812
rect 6788 11772 6794 11784
rect 7834 11772 7840 11784
rect 7892 11812 7898 11824
rect 7892 11784 7972 11812
rect 7892 11772 7898 11784
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 7006 11744 7012 11756
rect 6687 11716 7012 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7006 11704 7012 11716
rect 7064 11744 7070 11756
rect 7944 11753 7972 11784
rect 8478 11772 8484 11824
rect 8536 11812 8542 11824
rect 9876 11812 9904 11852
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 10008 11852 10425 11880
rect 10008 11840 10014 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 11514 11880 11520 11892
rect 10413 11843 10471 11849
rect 10888 11852 11520 11880
rect 10686 11812 10692 11824
rect 8536 11784 8694 11812
rect 9876 11784 10692 11812
rect 8536 11772 8542 11784
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7064 11716 7297 11744
rect 7064 11704 7070 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 9916 11716 10333 11744
rect 9916 11704 9922 11716
rect 10321 11713 10333 11716
rect 10367 11744 10379 11747
rect 10888 11744 10916 11852
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 13998 11880 14004 11892
rect 11756 11852 14004 11880
rect 11756 11840 11762 11852
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 14700 11852 15761 11880
rect 14700 11840 14706 11852
rect 15749 11849 15761 11852
rect 15795 11880 15807 11883
rect 16758 11880 16764 11892
rect 15795 11852 16764 11880
rect 15795 11849 15807 11852
rect 15749 11843 15807 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 18598 11880 18604 11892
rect 16868 11852 18604 11880
rect 11974 11812 11980 11824
rect 11935 11784 11980 11812
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 12434 11772 12440 11824
rect 12492 11772 12498 11824
rect 10367 11716 10916 11744
rect 10965 11747 11023 11753
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11422 11744 11428 11756
rect 11011 11716 11428 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 11698 11744 11704 11756
rect 11659 11716 11704 11744
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 14016 11753 14044 11840
rect 14277 11815 14335 11821
rect 14277 11781 14289 11815
rect 14323 11812 14335 11815
rect 14550 11812 14556 11824
rect 14323 11784 14556 11812
rect 14323 11781 14335 11784
rect 14277 11775 14335 11781
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 14734 11772 14740 11824
rect 14792 11772 14798 11824
rect 16868 11812 16896 11852
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 22094 11880 22100 11892
rect 19076 11852 22100 11880
rect 15580 11784 16896 11812
rect 17037 11815 17095 11821
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 5828 11648 6745 11676
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 11146 11676 11152 11688
rect 8251 11648 11152 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 11296 11648 13461 11676
rect 11296 11636 11302 11648
rect 13449 11645 13461 11648
rect 13495 11676 13507 11679
rect 15580 11676 15608 11784
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 17954 11812 17960 11824
rect 17083 11784 17960 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 19076 11821 19104 11852
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 24854 11880 24860 11892
rect 24815 11852 24860 11880
rect 24854 11840 24860 11852
rect 24912 11840 24918 11892
rect 19061 11815 19119 11821
rect 19061 11781 19073 11815
rect 19107 11781 19119 11815
rect 19061 11775 19119 11781
rect 20533 11815 20591 11821
rect 20533 11781 20545 11815
rect 20579 11812 20591 11815
rect 20622 11812 20628 11824
rect 20579 11784 20628 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 22189 11815 22247 11821
rect 22189 11812 22201 11815
rect 20772 11784 22201 11812
rect 20772 11772 20778 11784
rect 22189 11781 22201 11784
rect 22235 11781 22247 11815
rect 23106 11812 23112 11824
rect 23067 11784 23112 11812
rect 22189 11775 22247 11781
rect 23106 11772 23112 11784
rect 23164 11772 23170 11824
rect 24136 11784 25728 11812
rect 21542 11744 21548 11756
rect 21284 11716 21548 11744
rect 16942 11676 16948 11688
rect 13495 11648 15608 11676
rect 16903 11648 16948 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 17092 11648 17233 11676
rect 17092 11636 17098 11648
rect 17221 11645 17233 11648
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18279 11648 18981 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 20438 11676 20444 11688
rect 20351 11648 20444 11676
rect 18969 11639 19027 11645
rect 20438 11636 20444 11648
rect 20496 11676 20502 11688
rect 21284 11676 21312 11716
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 23566 11704 23572 11756
rect 23624 11744 23630 11756
rect 24026 11744 24032 11756
rect 23624 11716 24032 11744
rect 23624 11704 23630 11716
rect 24026 11704 24032 11716
rect 24084 11744 24090 11756
rect 24136 11753 24164 11784
rect 24121 11747 24179 11753
rect 24121 11744 24133 11747
rect 24084 11716 24133 11744
rect 24084 11704 24090 11716
rect 24121 11713 24133 11716
rect 24167 11713 24179 11747
rect 24762 11744 24768 11756
rect 24723 11716 24768 11744
rect 24121 11707 24179 11713
rect 24762 11704 24768 11716
rect 24820 11704 24826 11756
rect 25700 11753 25728 11784
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11713 25743 11747
rect 25685 11707 25743 11713
rect 29641 11747 29699 11753
rect 29641 11713 29653 11747
rect 29687 11744 29699 11747
rect 38102 11744 38108 11756
rect 29687 11716 38108 11744
rect 29687 11713 29699 11716
rect 29641 11707 29699 11713
rect 38102 11704 38108 11716
rect 38160 11704 38166 11756
rect 20496 11648 21312 11676
rect 21361 11679 21419 11685
rect 20496 11636 20502 11648
rect 21361 11645 21373 11679
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11676 22155 11679
rect 22186 11676 22192 11688
rect 22143 11648 22192 11676
rect 22143 11645 22155 11648
rect 22097 11639 22155 11645
rect 7650 11608 7656 11620
rect 5644 11580 7656 11608
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 10410 11608 10416 11620
rect 9600 11580 10416 11608
rect 5258 11540 5264 11552
rect 4172 11512 5264 11540
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5592 11512 6009 11540
rect 5592 11500 5598 11512
rect 5997 11509 6009 11512
rect 6043 11509 6055 11543
rect 5997 11503 6055 11509
rect 7377 11543 7435 11549
rect 7377 11509 7389 11543
rect 7423 11540 7435 11543
rect 9600 11540 9628 11580
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 17126 11608 17132 11620
rect 15672 11580 17132 11608
rect 7423 11512 9628 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 11057 11543 11115 11549
rect 9732 11512 9777 11540
rect 9732 11500 9738 11512
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 12526 11540 12532 11552
rect 11103 11512 12532 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 13446 11500 13452 11552
rect 13504 11540 13510 11552
rect 15672 11540 15700 11580
rect 17126 11568 17132 11580
rect 17184 11568 17190 11620
rect 19521 11611 19579 11617
rect 19521 11577 19533 11611
rect 19567 11577 19579 11611
rect 19521 11571 19579 11577
rect 13504 11512 15700 11540
rect 13504 11500 13510 11512
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 17034 11540 17040 11552
rect 15804 11512 17040 11540
rect 15804 11500 15810 11512
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 19536 11540 19564 11571
rect 21174 11568 21180 11620
rect 21232 11608 21238 11620
rect 21376 11608 21404 11639
rect 22186 11636 22192 11648
rect 22244 11676 22250 11688
rect 22244 11648 28994 11676
rect 22244 11636 22250 11648
rect 23106 11608 23112 11620
rect 21232 11580 23112 11608
rect 21232 11568 21238 11580
rect 23106 11568 23112 11580
rect 23164 11568 23170 11620
rect 21634 11540 21640 11552
rect 17276 11512 21640 11540
rect 17276 11500 17282 11512
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 21726 11500 21732 11552
rect 21784 11540 21790 11552
rect 22462 11540 22468 11552
rect 21784 11512 22468 11540
rect 21784 11500 21790 11512
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 22554 11500 22560 11552
rect 22612 11540 22618 11552
rect 24213 11543 24271 11549
rect 24213 11540 24225 11543
rect 22612 11512 24225 11540
rect 22612 11500 22618 11512
rect 24213 11509 24225 11512
rect 24259 11509 24271 11543
rect 24213 11503 24271 11509
rect 25501 11543 25559 11549
rect 25501 11509 25513 11543
rect 25547 11540 25559 11543
rect 26142 11540 26148 11552
rect 25547 11512 26148 11540
rect 25547 11509 25559 11512
rect 25501 11503 25559 11509
rect 26142 11500 26148 11512
rect 26200 11500 26206 11552
rect 28966 11540 28994 11648
rect 29733 11543 29791 11549
rect 29733 11540 29745 11543
rect 28966 11512 29745 11540
rect 29733 11509 29745 11512
rect 29779 11509 29791 11543
rect 29733 11503 29791 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 5718 11336 5724 11348
rect 2976 11308 5724 11336
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 2976 11118 3004 11308
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 6089 11339 6147 11345
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 6730 11336 6736 11348
rect 6135 11308 6736 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 6904 11339 6962 11345
rect 6904 11305 6916 11339
rect 6950 11336 6962 11339
rect 7558 11336 7564 11348
rect 6950 11308 7564 11336
rect 6950 11305 6962 11308
rect 6904 11299 6962 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 8389 11339 8447 11345
rect 7708 11308 8340 11336
rect 7708 11296 7714 11308
rect 8018 11228 8024 11280
rect 8076 11228 8082 11280
rect 8312 11268 8340 11308
rect 8389 11305 8401 11339
rect 8435 11336 8447 11339
rect 8662 11336 8668 11348
rect 8435 11308 8668 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9950 11336 9956 11348
rect 9911 11308 9956 11336
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 10376 11308 10609 11336
rect 10376 11296 10382 11308
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 10597 11299 10655 11305
rect 11256 11308 16160 11336
rect 9214 11268 9220 11280
rect 8312 11240 9220 11268
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 9309 11271 9367 11277
rect 9309 11237 9321 11271
rect 9355 11268 9367 11271
rect 11256 11268 11284 11308
rect 12894 11268 12900 11280
rect 9355 11240 11284 11268
rect 12855 11240 12900 11268
rect 9355 11237 9367 11240
rect 9309 11231 9367 11237
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 13633 11271 13691 11277
rect 13633 11237 13645 11271
rect 13679 11268 13691 11271
rect 13722 11268 13728 11280
rect 13679 11240 13728 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 3510 11200 3516 11212
rect 3375 11172 3516 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 4304 11172 4353 11200
rect 4304 11160 4310 11172
rect 4341 11169 4353 11172
rect 4387 11200 4399 11203
rect 4614 11200 4620 11212
rect 4387 11172 4620 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5810 11200 5816 11212
rect 5316 11172 5816 11200
rect 5316 11160 5322 11172
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6641 11203 6699 11209
rect 6641 11169 6653 11203
rect 6687 11200 6699 11203
rect 8036 11200 8064 11228
rect 6687 11172 8064 11200
rect 6687 11169 6699 11172
rect 6641 11163 6699 11169
rect 8386 11160 8392 11212
rect 8444 11200 8450 11212
rect 8938 11200 8944 11212
rect 8444 11172 8944 11200
rect 8444 11160 8450 11172
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9030 11160 9036 11212
rect 9088 11200 9094 11212
rect 9088 11172 10088 11200
rect 9088 11160 9094 11172
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 8260 11104 9229 11132
rect 8260 11092 8266 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 9861 11135 9919 11141
rect 9861 11132 9873 11135
rect 9732 11104 9873 11132
rect 9732 11092 9738 11104
rect 9861 11101 9873 11104
rect 9907 11101 9919 11135
rect 10060 11132 10088 11172
rect 11974 11160 11980 11212
rect 12032 11200 12038 11212
rect 13446 11200 13452 11212
rect 12032 11172 13452 11200
rect 12032 11160 12038 11172
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 14608 11172 16037 11200
rect 14608 11160 14614 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 10060 11104 10517 11132
rect 9861 11095 9919 11101
rect 10505 11101 10517 11104
rect 10551 11132 10563 11135
rect 10594 11132 10600 11144
rect 10551 11104 10600 11132
rect 10551 11101 10563 11104
rect 10505 11095 10563 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11146 11132 11152 11144
rect 11107 11104 11152 11132
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 12952 11104 13553 11132
rect 12952 11092 12958 11104
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 14056 11104 14289 11132
rect 14056 11092 14062 11104
rect 14277 11101 14289 11104
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 1026 11024 1032 11076
rect 1084 11064 1090 11076
rect 1302 11064 1308 11076
rect 1084 11036 1308 11064
rect 1084 11024 1090 11036
rect 1302 11024 1308 11036
rect 1360 11064 1366 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1360 11036 1869 11064
rect 1360 11024 1366 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 4614 11064 4620 11076
rect 1857 11027 1915 11033
rect 3252 11036 3464 11064
rect 4575 11036 4620 11064
rect 1762 10956 1768 11008
rect 1820 10996 1826 11008
rect 3252 10996 3280 11036
rect 1820 10968 3280 10996
rect 3436 10996 3464 11036
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 7190 11064 7196 11076
rect 5842 11036 7196 11064
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7374 11024 7380 11076
rect 7432 11024 7438 11076
rect 9232 11036 10088 11064
rect 9232 10996 9260 11036
rect 3436 10968 9260 10996
rect 10060 10996 10088 11036
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 11388 11036 11437 11064
rect 11388 11024 11394 11036
rect 11425 11033 11437 11036
rect 11471 11033 11483 11067
rect 11425 11027 11483 11033
rect 11882 11024 11888 11076
rect 11940 11024 11946 11076
rect 13722 11024 13728 11076
rect 13780 11064 13786 11076
rect 14550 11064 14556 11076
rect 13780 11036 14412 11064
rect 14511 11036 14556 11064
rect 13780 11024 13786 11036
rect 12434 10996 12440 11008
rect 10060 10968 12440 10996
rect 1820 10956 1826 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 14384 10996 14412 11036
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 16132 11064 16160 11308
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 21726 11336 21732 11348
rect 18012 11308 21732 11336
rect 18012 11296 18018 11308
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 24762 11336 24768 11348
rect 21836 11308 24768 11336
rect 16298 11228 16304 11280
rect 16356 11268 16362 11280
rect 16356 11240 16712 11268
rect 16356 11228 16362 11240
rect 16574 11200 16580 11212
rect 16535 11172 16580 11200
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 16684 11200 16712 11240
rect 17034 11228 17040 11280
rect 17092 11268 17098 11280
rect 17092 11240 19472 11268
rect 17092 11228 17098 11240
rect 18233 11203 18291 11209
rect 18233 11200 18245 11203
rect 16684 11172 18245 11200
rect 18233 11169 18245 11172
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11132 18107 11135
rect 18414 11132 18420 11144
rect 18095 11104 18420 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 19444 11141 19472 11240
rect 20438 11228 20444 11280
rect 20496 11268 20502 11280
rect 21836 11268 21864 11308
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 38102 11336 38108 11348
rect 38063 11308 38108 11336
rect 38102 11296 38108 11308
rect 38160 11296 38166 11348
rect 20496 11240 21864 11268
rect 20496 11228 20502 11240
rect 21910 11228 21916 11280
rect 21968 11268 21974 11280
rect 26878 11268 26884 11280
rect 21968 11240 26884 11268
rect 21968 11228 21974 11240
rect 26878 11228 26884 11240
rect 26936 11228 26942 11280
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11200 20223 11203
rect 22186 11200 22192 11212
rect 20211 11172 22192 11200
rect 20211 11169 20223 11172
rect 20165 11163 20223 11169
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 23290 11132 23296 11144
rect 19429 11095 19487 11101
rect 21008 11104 21312 11132
rect 23251 11104 23296 11132
rect 21008 11076 21036 11104
rect 16669 11067 16727 11073
rect 16669 11064 16681 11067
rect 14660 11036 15042 11064
rect 16132 11036 16681 11064
rect 14660 10996 14688 11036
rect 16669 11033 16681 11036
rect 16715 11033 16727 11067
rect 16669 11027 16727 11033
rect 17218 11024 17224 11076
rect 17276 11064 17282 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17276 11036 17601 11064
rect 17276 11024 17282 11036
rect 17589 11033 17601 11036
rect 17635 11033 17647 11067
rect 17589 11027 17647 11033
rect 19521 11067 19579 11073
rect 19521 11033 19533 11067
rect 19567 11064 19579 11067
rect 20257 11067 20315 11073
rect 19567 11036 20116 11064
rect 19567 11033 19579 11036
rect 19521 11027 19579 11033
rect 14384 10968 14688 10996
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 19334 10996 19340 11008
rect 14884 10968 19340 10996
rect 14884 10956 14890 10968
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 20088 10996 20116 11036
rect 20257 11033 20269 11067
rect 20303 11033 20315 11067
rect 20257 11027 20315 11033
rect 20272 10996 20300 11027
rect 20622 11024 20628 11076
rect 20680 11064 20686 11076
rect 20990 11064 20996 11076
rect 20680 11036 20996 11064
rect 20680 11024 20686 11036
rect 20990 11024 20996 11036
rect 21048 11024 21054 11076
rect 21082 11024 21088 11076
rect 21140 11064 21146 11076
rect 21177 11067 21235 11073
rect 21177 11064 21189 11067
rect 21140 11036 21189 11064
rect 21140 11024 21146 11036
rect 21177 11033 21189 11036
rect 21223 11033 21235 11067
rect 21284 11064 21312 11104
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 26142 11132 26148 11144
rect 26103 11104 26148 11132
rect 24765 11095 24823 11101
rect 21821 11067 21879 11073
rect 21821 11064 21833 11067
rect 21284 11036 21833 11064
rect 21177 11027 21235 11033
rect 21821 11033 21833 11036
rect 21867 11033 21879 11067
rect 21821 11027 21879 11033
rect 21910 11024 21916 11076
rect 21968 11064 21974 11076
rect 22830 11064 22836 11076
rect 21968 11036 22013 11064
rect 22791 11036 22836 11064
rect 21968 11024 21974 11036
rect 22830 11024 22836 11036
rect 22888 11024 22894 11076
rect 23106 11024 23112 11076
rect 23164 11064 23170 11076
rect 24780 11064 24808 11095
rect 26142 11092 26148 11104
rect 26200 11092 26206 11144
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 23164 11036 24808 11064
rect 23164 11024 23170 11036
rect 20088 10968 20300 10996
rect 20530 10956 20536 11008
rect 20588 10996 20594 11008
rect 23385 10999 23443 11005
rect 23385 10996 23397 10999
rect 20588 10968 23397 10996
rect 20588 10956 20594 10968
rect 23385 10965 23397 10968
rect 23431 10965 23443 10999
rect 23385 10959 23443 10965
rect 24581 10999 24639 11005
rect 24581 10965 24593 10999
rect 24627 10996 24639 10999
rect 24762 10996 24768 11008
rect 24627 10968 24768 10996
rect 24627 10965 24639 10968
rect 24581 10959 24639 10965
rect 24762 10956 24768 10968
rect 24820 10956 24826 11008
rect 25958 10996 25964 11008
rect 25919 10968 25964 10996
rect 25958 10956 25964 10968
rect 26016 10956 26022 11008
rect 26602 10996 26608 11008
rect 26563 10968 26608 10996
rect 26602 10956 26608 10968
rect 26660 10956 26666 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1762 10792 1768 10804
rect 1723 10764 1768 10792
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2314 10792 2320 10804
rect 2275 10764 2320 10792
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 2498 10752 2504 10804
rect 2556 10792 2562 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 2556 10764 3065 10792
rect 2556 10752 2562 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3384 10764 3709 10792
rect 3384 10752 3390 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 3697 10755 3755 10761
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10792 6055 10795
rect 6454 10792 6460 10804
rect 6043 10764 6460 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6454 10752 6460 10764
rect 6512 10792 6518 10804
rect 6638 10792 6644 10804
rect 6512 10764 6644 10792
rect 6512 10752 6518 10764
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7285 10795 7343 10801
rect 7285 10761 7297 10795
rect 7331 10792 7343 10795
rect 11057 10795 11115 10801
rect 7331 10764 10732 10792
rect 7331 10761 7343 10764
rect 7285 10755 7343 10761
rect 934 10684 940 10736
rect 992 10724 998 10736
rect 992 10696 2544 10724
rect 992 10684 998 10696
rect 2516 10665 2544 10696
rect 3418 10684 3424 10736
rect 3476 10724 3482 10736
rect 4525 10727 4583 10733
rect 4525 10724 4537 10727
rect 3476 10696 4537 10724
rect 3476 10684 3482 10696
rect 4525 10693 4537 10696
rect 4571 10693 4583 10727
rect 6822 10724 6828 10736
rect 5750 10696 6828 10724
rect 4525 10687 4583 10693
rect 6822 10684 6828 10696
rect 6880 10684 6886 10736
rect 7742 10724 7748 10736
rect 7116 10696 7748 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3050 10656 3056 10668
rect 3007 10628 3056 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 1688 10588 1716 10619
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10625 3663 10659
rect 4246 10656 4252 10668
rect 4207 10628 4252 10656
rect 3605 10619 3663 10625
rect 3620 10588 3648 10619
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 7116 10656 7144 10696
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 8018 10724 8024 10736
rect 7852 10696 8024 10724
rect 6595 10628 7144 10656
rect 7193 10659 7251 10665
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7282 10656 7288 10668
rect 7239 10628 7288 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7852 10665 7880 10696
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 8113 10727 8171 10733
rect 8113 10693 8125 10727
rect 8159 10724 8171 10727
rect 8386 10724 8392 10736
rect 8159 10696 8392 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 8386 10684 8392 10696
rect 8444 10684 8450 10736
rect 10594 10724 10600 10736
rect 9338 10696 10600 10724
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 10704 10724 10732 10764
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11882 10792 11888 10804
rect 11103 10764 11888 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12158 10752 12164 10804
rect 12216 10792 12222 10804
rect 12216 10764 15792 10792
rect 12216 10752 12222 10764
rect 12250 10724 12256 10736
rect 10704 10696 12256 10724
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 13262 10684 13268 10736
rect 13320 10724 13326 10736
rect 14277 10727 14335 10733
rect 14277 10724 14289 10727
rect 13320 10696 14289 10724
rect 13320 10684 13326 10696
rect 14277 10693 14289 10696
rect 14323 10693 14335 10727
rect 15654 10724 15660 10736
rect 15502 10696 15660 10724
rect 14277 10687 14335 10693
rect 15654 10684 15660 10696
rect 15712 10684 15718 10736
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 10134 10656 10140 10668
rect 7837 10619 7895 10625
rect 9508 10628 10140 10656
rect 9508 10588 9536 10628
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10284 10628 10333 10656
rect 10284 10616 10290 10628
rect 10321 10625 10333 10628
rect 10367 10656 10379 10659
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10367 10628 10977 10656
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 10965 10625 10977 10628
rect 11011 10656 11023 10659
rect 11330 10656 11336 10668
rect 11011 10628 11336 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 13110 10628 13860 10656
rect 1688 10560 2774 10588
rect 3620 10560 9536 10588
rect 9585 10591 9643 10597
rect 2746 10520 2774 10560
rect 9585 10557 9597 10591
rect 9631 10588 9643 10591
rect 11054 10588 11060 10600
rect 9631 10560 11060 10588
rect 9631 10557 9643 10560
rect 9585 10551 9643 10557
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 11698 10588 11704 10600
rect 11659 10560 11704 10588
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10588 12035 10591
rect 12066 10588 12072 10600
rect 12023 10560 12072 10588
rect 12023 10557 12035 10560
rect 11977 10551 12035 10557
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 12400 10560 13461 10588
rect 12400 10548 12406 10560
rect 13449 10557 13461 10560
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 3786 10520 3792 10532
rect 2746 10492 3792 10520
rect 3786 10480 3792 10492
rect 3844 10480 3850 10532
rect 7834 10520 7840 10532
rect 6472 10492 7840 10520
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 6472 10452 6500 10492
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 10413 10523 10471 10529
rect 10413 10489 10425 10523
rect 10459 10520 10471 10523
rect 10459 10492 11468 10520
rect 10459 10489 10471 10492
rect 10413 10483 10471 10489
rect 6638 10452 6644 10464
rect 5316 10424 6500 10452
rect 6599 10424 6644 10452
rect 5316 10412 5322 10424
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7282 10452 7288 10464
rect 7156 10424 7288 10452
rect 7156 10412 7162 10424
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 9674 10452 9680 10464
rect 7524 10424 9680 10452
rect 7524 10412 7530 10424
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10778 10452 10784 10464
rect 10560 10424 10784 10452
rect 10560 10412 10566 10424
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11440 10452 11468 10492
rect 13722 10452 13728 10464
rect 11440 10424 13728 10452
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 13832 10452 13860 10628
rect 13998 10588 14004 10600
rect 13959 10560 14004 10588
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 14826 10588 14832 10600
rect 14332 10560 14832 10588
rect 14332 10548 14338 10560
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 14826 10452 14832 10464
rect 13832 10424 14832 10452
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 15764 10461 15792 10764
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 23569 10795 23627 10801
rect 23569 10792 23581 10795
rect 18932 10764 23581 10792
rect 18932 10752 18938 10764
rect 23569 10761 23581 10764
rect 23615 10761 23627 10795
rect 24118 10792 24124 10804
rect 24079 10764 24124 10792
rect 23569 10755 23627 10761
rect 24118 10752 24124 10764
rect 24176 10752 24182 10804
rect 17494 10724 17500 10736
rect 16868 10696 17500 10724
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 16868 10665 16896 10696
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 18506 10724 18512 10736
rect 18467 10696 18512 10724
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 19426 10724 19432 10736
rect 19387 10696 19432 10724
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 20257 10727 20315 10733
rect 20257 10693 20269 10727
rect 20303 10724 20315 10727
rect 20806 10724 20812 10736
rect 20303 10696 20812 10724
rect 20303 10693 20315 10696
rect 20257 10687 20315 10693
rect 20806 10684 20812 10696
rect 20864 10684 20870 10736
rect 21174 10724 21180 10736
rect 21135 10696 21180 10724
rect 21174 10684 21180 10696
rect 21232 10684 21238 10736
rect 21266 10684 21272 10736
rect 21324 10724 21330 10736
rect 22002 10724 22008 10736
rect 21324 10696 22008 10724
rect 21324 10684 21330 10696
rect 22002 10684 22008 10696
rect 22060 10724 22066 10736
rect 25866 10724 25872 10736
rect 22060 10696 23520 10724
rect 22060 10684 22066 10696
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16816 10628 16865 10656
rect 16816 10616 16822 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17310 10656 17316 10668
rect 17083 10628 17316 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 21542 10616 21548 10668
rect 21600 10656 21606 10668
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 21600 10628 22385 10656
rect 21600 10616 21606 10628
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22554 10656 22560 10668
rect 22515 10628 22560 10656
rect 22373 10619 22431 10625
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 23492 10665 23520 10696
rect 23952 10696 25872 10724
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10625 23535 10659
rect 23477 10619 23535 10625
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 17000 10560 18429 10588
rect 17000 10548 17006 10560
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 18506 10548 18512 10600
rect 18564 10588 18570 10600
rect 18874 10588 18880 10600
rect 18564 10560 18880 10588
rect 18564 10548 18570 10560
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 19058 10548 19064 10600
rect 19116 10588 19122 10600
rect 19978 10588 19984 10600
rect 19116 10560 19984 10588
rect 19116 10548 19122 10560
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 21082 10588 21088 10600
rect 20211 10560 21088 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 21082 10548 21088 10560
rect 21140 10548 21146 10600
rect 22094 10548 22100 10600
rect 22152 10588 22158 10600
rect 23952 10588 23980 10696
rect 25866 10684 25872 10696
rect 25924 10724 25930 10736
rect 29365 10727 29423 10733
rect 29365 10724 29377 10727
rect 25924 10696 29377 10724
rect 25924 10684 25930 10696
rect 29365 10693 29377 10696
rect 29411 10693 29423 10727
rect 29365 10687 29423 10693
rect 25958 10656 25964 10668
rect 25919 10628 25964 10656
rect 25958 10616 25964 10628
rect 26016 10616 26022 10668
rect 29273 10659 29331 10665
rect 29273 10625 29285 10659
rect 29319 10625 29331 10659
rect 29273 10619 29331 10625
rect 30837 10659 30895 10665
rect 30837 10625 30849 10659
rect 30883 10656 30895 10659
rect 33042 10656 33048 10668
rect 30883 10628 33048 10656
rect 30883 10625 30895 10628
rect 30837 10619 30895 10625
rect 22152 10560 23980 10588
rect 22152 10548 22158 10560
rect 24210 10548 24216 10600
rect 24268 10588 24274 10600
rect 24765 10591 24823 10597
rect 24765 10588 24777 10591
rect 24268 10560 24777 10588
rect 24268 10548 24274 10560
rect 24765 10557 24777 10560
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 25777 10591 25835 10597
rect 25777 10557 25789 10591
rect 25823 10588 25835 10591
rect 26602 10588 26608 10600
rect 25823 10560 26608 10588
rect 25823 10557 25835 10560
rect 25777 10551 25835 10557
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 29288 10588 29316 10619
rect 33042 10616 33048 10628
rect 33100 10616 33106 10668
rect 38102 10588 38108 10600
rect 29288 10560 38108 10588
rect 38102 10548 38108 10560
rect 38160 10548 38166 10600
rect 16482 10480 16488 10532
rect 16540 10520 16546 10532
rect 17221 10523 17279 10529
rect 17221 10520 17233 10523
rect 16540 10492 17233 10520
rect 16540 10480 16546 10492
rect 17221 10489 17233 10492
rect 17267 10489 17279 10523
rect 23106 10520 23112 10532
rect 17221 10483 17279 10489
rect 17328 10492 23112 10520
rect 15749 10455 15807 10461
rect 15749 10421 15761 10455
rect 15795 10452 15807 10455
rect 17328 10452 17356 10492
rect 23106 10480 23112 10492
rect 23164 10480 23170 10532
rect 15795 10424 17356 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 20990 10452 20996 10464
rect 17552 10424 20996 10452
rect 17552 10412 17558 10424
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 21174 10412 21180 10464
rect 21232 10452 21238 10464
rect 22922 10452 22928 10464
rect 21232 10424 22928 10452
rect 21232 10412 21238 10424
rect 22922 10412 22928 10424
rect 22980 10412 22986 10464
rect 23017 10455 23075 10461
rect 23017 10421 23029 10455
rect 23063 10452 23075 10455
rect 24486 10452 24492 10464
rect 23063 10424 24492 10452
rect 23063 10421 23075 10424
rect 23017 10415 23075 10421
rect 24486 10412 24492 10424
rect 24544 10452 24550 10464
rect 26145 10455 26203 10461
rect 26145 10452 26157 10455
rect 24544 10424 26157 10452
rect 24544 10412 24550 10424
rect 26145 10421 26157 10424
rect 26191 10421 26203 10455
rect 30926 10452 30932 10464
rect 30887 10424 30932 10452
rect 26145 10415 26203 10421
rect 30926 10412 30932 10424
rect 30984 10412 30990 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3016 10220 3433 10248
rect 3016 10208 3022 10220
rect 3421 10217 3433 10220
rect 3467 10248 3479 10251
rect 5626 10248 5632 10260
rect 3467 10220 5632 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 6638 10208 6644 10260
rect 6696 10248 6702 10260
rect 16390 10248 16396 10260
rect 6696 10220 16396 10248
rect 6696 10208 6702 10220
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16574 10248 16580 10260
rect 16535 10220 16580 10248
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 19702 10248 19708 10260
rect 18288 10220 19708 10248
rect 18288 10208 18294 10220
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 22278 10208 22284 10260
rect 22336 10248 22342 10260
rect 22465 10251 22523 10257
rect 22465 10248 22477 10251
rect 22336 10220 22477 10248
rect 22336 10208 22342 10220
rect 22465 10217 22477 10220
rect 22511 10217 22523 10251
rect 22465 10211 22523 10217
rect 22922 10208 22928 10260
rect 22980 10248 22986 10260
rect 25317 10251 25375 10257
rect 25317 10248 25329 10251
rect 22980 10220 25329 10248
rect 22980 10208 22986 10220
rect 25317 10217 25329 10220
rect 25363 10217 25375 10251
rect 25317 10211 25375 10217
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 11330 10180 11336 10192
rect 8444 10152 11336 10180
rect 8444 10140 8450 10152
rect 11330 10140 11336 10152
rect 11388 10180 11394 10192
rect 11882 10180 11888 10192
rect 11388 10152 11888 10180
rect 11388 10140 11394 10152
rect 11882 10140 11888 10152
rect 11940 10140 11946 10192
rect 13446 10140 13452 10192
rect 13504 10180 13510 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 13504 10152 13645 10180
rect 13504 10140 13510 10152
rect 13633 10149 13645 10152
rect 13679 10149 13691 10183
rect 13633 10143 13691 10149
rect 15838 10140 15844 10192
rect 15896 10180 15902 10192
rect 16850 10180 16856 10192
rect 15896 10152 16856 10180
rect 15896 10140 15902 10152
rect 16850 10140 16856 10152
rect 16908 10180 16914 10192
rect 19058 10180 19064 10192
rect 16908 10152 19064 10180
rect 16908 10140 16914 10152
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 19426 10180 19432 10192
rect 19306 10152 19432 10180
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2590 10112 2596 10124
rect 1719 10084 2596 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2590 10072 2596 10084
rect 2648 10112 2654 10124
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 2648 10084 3985 10112
rect 2648 10072 2654 10084
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 6822 10112 6828 10124
rect 5960 10084 6040 10112
rect 6783 10084 6828 10112
rect 5960 10072 5966 10084
rect 6012 10053 6040 10084
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7466 10112 7472 10124
rect 7147 10084 7472 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7466 10072 7472 10084
rect 7524 10112 7530 10124
rect 7650 10112 7656 10124
rect 7524 10084 7656 10112
rect 7524 10072 7530 10084
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 11054 10112 11060 10124
rect 7800 10084 11060 10112
rect 7800 10072 7806 10084
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10112 14703 10115
rect 14918 10112 14924 10124
rect 14691 10084 14924 10112
rect 14691 10081 14703 10084
rect 14645 10075 14703 10081
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 15562 10112 15568 10124
rect 15523 10084 15568 10112
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10112 17371 10115
rect 17402 10112 17408 10124
rect 17359 10084 17408 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 18690 10112 18696 10124
rect 18603 10084 18696 10112
rect 18690 10072 18696 10084
rect 18748 10112 18754 10124
rect 19306 10112 19334 10152
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 20073 10183 20131 10189
rect 20073 10149 20085 10183
rect 20119 10180 20131 10183
rect 20254 10180 20260 10192
rect 20119 10152 20260 10180
rect 20119 10149 20131 10152
rect 20073 10143 20131 10149
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 18748 10084 19334 10112
rect 19522 10115 19580 10121
rect 18748 10072 18754 10084
rect 19522 10081 19534 10115
rect 19568 10112 19580 10115
rect 19886 10112 19892 10124
rect 19568 10084 19892 10112
rect 19568 10081 19580 10084
rect 19522 10075 19580 10081
rect 19886 10072 19892 10084
rect 19944 10072 19950 10124
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 21634 10112 21640 10124
rect 20036 10084 21640 10112
rect 20036 10072 20042 10084
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 23201 10115 23259 10121
rect 23201 10081 23213 10115
rect 23247 10112 23259 10115
rect 24210 10112 24216 10124
rect 23247 10084 24216 10112
rect 23247 10081 23259 10084
rect 23201 10075 23259 10081
rect 24210 10072 24216 10084
rect 24268 10072 24274 10124
rect 25240 10084 33180 10112
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10044 6055 10047
rect 6638 10044 6644 10056
rect 6043 10016 6644 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16206 10044 16212 10056
rect 16163 10016 16212 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 1946 9976 1952 9988
rect 1907 9948 1952 9976
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 3174 9948 3464 9976
rect 3436 9908 3464 9948
rect 3510 9936 3516 9988
rect 3568 9976 3574 9988
rect 4249 9979 4307 9985
rect 4249 9976 4261 9979
rect 3568 9948 4261 9976
rect 3568 9936 3574 9948
rect 4249 9945 4261 9948
rect 4295 9945 4307 9979
rect 5902 9976 5908 9988
rect 5474 9948 5908 9976
rect 4249 9939 4307 9945
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 9125 9979 9183 9985
rect 9125 9976 9137 9979
rect 6012 9948 7590 9976
rect 8404 9948 9137 9976
rect 5074 9908 5080 9920
rect 3436 9880 5080 9908
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5258 9868 5264 9920
rect 5316 9908 5322 9920
rect 6012 9908 6040 9948
rect 5316 9880 6040 9908
rect 5316 9868 5322 9880
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 8404 9908 8432 9948
rect 9125 9945 9137 9948
rect 9171 9945 9183 9979
rect 9125 9939 9183 9945
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 11900 9976 11928 10007
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10044 16359 10047
rect 16666 10044 16672 10056
rect 16347 10016 16672 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 18414 10044 18420 10056
rect 18375 10016 18420 10044
rect 18414 10004 18420 10016
rect 18472 10044 18478 10056
rect 19150 10044 19156 10056
rect 18472 10016 19156 10044
rect 18472 10004 18478 10016
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 24762 10044 24768 10056
rect 24723 10016 24768 10044
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 25240 10053 25268 10084
rect 25225 10047 25283 10053
rect 25225 10013 25237 10047
rect 25271 10013 25283 10047
rect 26050 10044 26056 10056
rect 26011 10016 26056 10044
rect 25225 10007 25283 10013
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 33152 9988 33180 10084
rect 34514 10072 34520 10124
rect 34572 10112 34578 10124
rect 37737 10115 37795 10121
rect 37737 10112 37749 10115
rect 34572 10084 37749 10112
rect 34572 10072 34578 10084
rect 37737 10081 37749 10084
rect 37783 10081 37795 10115
rect 37737 10075 37795 10081
rect 37182 10004 37188 10056
rect 37240 10044 37246 10056
rect 37461 10047 37519 10053
rect 37461 10044 37473 10047
rect 37240 10016 37473 10044
rect 37240 10004 37246 10016
rect 37461 10013 37473 10016
rect 37507 10013 37519 10047
rect 37461 10007 37519 10013
rect 12158 9976 12164 9988
rect 11204 9948 11928 9976
rect 12119 9948 12164 9976
rect 11204 9936 11210 9948
rect 12158 9936 12164 9948
rect 12216 9936 12222 9988
rect 12802 9936 12808 9988
rect 12860 9936 12866 9988
rect 13722 9936 13728 9988
rect 13780 9976 13786 9988
rect 14737 9979 14795 9985
rect 14737 9976 14749 9979
rect 13780 9948 14749 9976
rect 13780 9936 13786 9948
rect 14737 9945 14749 9948
rect 14783 9945 14795 9979
rect 14737 9939 14795 9945
rect 16390 9936 16396 9988
rect 16448 9976 16454 9988
rect 17405 9979 17463 9985
rect 17405 9976 17417 9979
rect 16448 9948 17417 9976
rect 16448 9936 16454 9948
rect 17405 9945 17417 9948
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 17957 9979 18015 9985
rect 17957 9945 17969 9979
rect 18003 9976 18015 9979
rect 18598 9976 18604 9988
rect 18003 9948 18604 9976
rect 18003 9945 18015 9948
rect 17957 9939 18015 9945
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 19518 9976 19524 9988
rect 19306 9948 19524 9976
rect 6144 9880 8432 9908
rect 6144 9868 6150 9880
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8536 9880 8585 9908
rect 8536 9868 8542 9880
rect 8573 9877 8585 9880
rect 8619 9908 8631 9911
rect 9674 9908 9680 9920
rect 8619 9880 9680 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 10413 9911 10471 9917
rect 10413 9908 10425 9911
rect 9824 9880 10425 9908
rect 9824 9868 9830 9880
rect 10413 9877 10425 9880
rect 10459 9877 10471 9911
rect 10413 9871 10471 9877
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 13078 9908 13084 9920
rect 10560 9880 13084 9908
rect 10560 9868 10566 9880
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 15930 9868 15936 9920
rect 15988 9908 15994 9920
rect 19306 9908 19334 9948
rect 19518 9936 19524 9948
rect 19576 9936 19582 9988
rect 19613 9979 19671 9985
rect 19613 9945 19625 9979
rect 19659 9976 19671 9979
rect 19659 9948 19840 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 15988 9880 19334 9908
rect 19812 9908 19840 9948
rect 19886 9936 19892 9988
rect 19944 9976 19950 9988
rect 21177 9979 21235 9985
rect 21177 9976 21189 9979
rect 19944 9948 21189 9976
rect 19944 9936 19950 9948
rect 21177 9945 21189 9948
rect 21223 9945 21235 9979
rect 21177 9939 21235 9945
rect 21269 9979 21327 9985
rect 21269 9945 21281 9979
rect 21315 9945 21327 9979
rect 21818 9976 21824 9988
rect 21779 9948 21824 9976
rect 21269 9939 21327 9945
rect 20530 9908 20536 9920
rect 19812 9880 20536 9908
rect 15988 9868 15994 9880
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 21284 9908 21312 9939
rect 21818 9936 21824 9948
rect 21876 9936 21882 9988
rect 22094 9936 22100 9988
rect 22152 9976 22158 9988
rect 22373 9979 22431 9985
rect 22373 9976 22385 9979
rect 22152 9948 22385 9976
rect 22152 9936 22158 9948
rect 22373 9945 22385 9948
rect 22419 9945 22431 9979
rect 22373 9939 22431 9945
rect 23293 9979 23351 9985
rect 23293 9945 23305 9979
rect 23339 9976 23351 9979
rect 23842 9976 23848 9988
rect 23339 9948 23520 9976
rect 23755 9948 23848 9976
rect 23339 9945 23351 9948
rect 23293 9939 23351 9945
rect 22738 9908 22744 9920
rect 21284 9880 22744 9908
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 23492 9908 23520 9948
rect 23842 9936 23848 9948
rect 23900 9976 23906 9988
rect 28258 9976 28264 9988
rect 23900 9948 28264 9976
rect 23900 9936 23906 9948
rect 28258 9936 28264 9948
rect 28316 9936 28322 9988
rect 33134 9936 33140 9988
rect 33192 9976 33198 9988
rect 34422 9976 34428 9988
rect 33192 9948 34428 9976
rect 33192 9936 33198 9948
rect 34422 9936 34428 9948
rect 34480 9936 34486 9988
rect 24581 9911 24639 9917
rect 24581 9908 24593 9911
rect 23492 9880 24593 9908
rect 24581 9877 24593 9880
rect 24627 9877 24639 9911
rect 24581 9871 24639 9877
rect 25869 9911 25927 9917
rect 25869 9877 25881 9911
rect 25915 9908 25927 9911
rect 25958 9908 25964 9920
rect 25915 9880 25964 9908
rect 25915 9877 25927 9880
rect 25869 9871 25927 9877
rect 25958 9868 25964 9880
rect 26016 9868 26022 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 10502 9704 10508 9716
rect 5960 9676 10508 9704
rect 5960 9664 5966 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 17402 9704 17408 9716
rect 15252 9676 17408 9704
rect 15252 9664 15258 9676
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 17954 9704 17960 9716
rect 17512 9676 17960 9704
rect 3510 9636 3516 9648
rect 3082 9608 3516 9636
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 8018 9636 8024 9648
rect 5750 9608 8024 9636
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 9582 9636 9588 9648
rect 8970 9608 9588 9636
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 13446 9636 13452 9648
rect 13386 9608 13452 9636
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 14182 9596 14188 9648
rect 14240 9636 14246 9648
rect 14369 9639 14427 9645
rect 14369 9636 14381 9639
rect 14240 9608 14381 9636
rect 14240 9596 14246 9608
rect 14369 9605 14381 9608
rect 14415 9605 14427 9639
rect 16022 9636 16028 9648
rect 14369 9599 14427 9605
rect 15856 9608 16028 9636
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 6546 9568 6552 9580
rect 5960 9540 6552 9568
rect 5960 9528 5966 9540
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 8956 9540 9720 9568
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 1857 9503 1915 9509
rect 1627 9472 1716 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 1688 9364 1716 9472
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2498 9500 2504 9512
rect 1903 9472 2504 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 3252 9472 4261 9500
rect 2222 9364 2228 9376
rect 1688 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9364 2286 9376
rect 2590 9364 2596 9376
rect 2280 9336 2596 9364
rect 2280 9324 2286 9336
rect 2590 9324 2596 9336
rect 2648 9364 2654 9376
rect 3252 9364 3280 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 5534 9500 5540 9512
rect 4571 9472 5540 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 2648 9336 3280 9364
rect 3329 9367 3387 9373
rect 2648 9324 2654 9336
rect 3329 9333 3341 9367
rect 3375 9364 3387 9367
rect 3418 9364 3424 9376
rect 3375 9336 3424 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 3418 9324 3424 9336
rect 3476 9364 3482 9376
rect 3878 9364 3884 9376
rect 3476 9336 3884 9364
rect 3476 9324 3482 9336
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 4264 9364 4292 9463
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 5994 9500 6000 9512
rect 5955 9472 6000 9500
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6546 9432 6552 9444
rect 6507 9404 6552 9432
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 4706 9364 4712 9376
rect 4264 9336 4712 9364
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 5166 9324 5172 9376
rect 5224 9364 5230 9376
rect 6748 9364 6776 9531
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7466 9500 7472 9512
rect 6972 9472 7472 9500
rect 6972 9460 6978 9472
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 7834 9500 7840 9512
rect 7791 9472 7840 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8956 9500 8984 9540
rect 8168 9472 8984 9500
rect 9493 9503 9551 9509
rect 8168 9460 8174 9472
rect 9493 9469 9505 9503
rect 9539 9469 9551 9503
rect 9692 9500 9720 9540
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9824 9540 9965 9568
rect 9824 9528 9830 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10560 9540 10701 9568
rect 10560 9528 10566 9540
rect 10689 9537 10701 9540
rect 10735 9568 10747 9571
rect 11146 9568 11152 9580
rect 10735 9540 11152 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 15856 9577 15884 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17512 9636 17540 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 20346 9704 20352 9716
rect 18064 9676 20352 9704
rect 17083 9608 17540 9636
rect 17589 9639 17647 9645
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17589 9605 17601 9639
rect 17635 9636 17647 9639
rect 17770 9636 17776 9648
rect 17635 9608 17776 9636
rect 17635 9605 17647 9608
rect 17589 9599 17647 9605
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 18064 9636 18092 9676
rect 20346 9664 20352 9676
rect 20404 9664 20410 9716
rect 21082 9664 21088 9716
rect 21140 9704 21146 9716
rect 30926 9704 30932 9716
rect 21140 9676 30932 9704
rect 21140 9664 21146 9676
rect 30926 9664 30932 9676
rect 30984 9664 30990 9716
rect 17880 9608 18092 9636
rect 18601 9639 18659 9645
rect 15841 9571 15899 9577
rect 13372 9540 15240 9568
rect 11790 9500 11796 9512
rect 9692 9472 11796 9500
rect 9493 9463 9551 9469
rect 5224 9336 6776 9364
rect 5224 9324 5230 9336
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 9508 9364 9536 9463
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9469 11943 9503
rect 12158 9500 12164 9512
rect 12071 9472 12164 9500
rect 11885 9463 11943 9469
rect 10410 9392 10416 9444
rect 10468 9432 10474 9444
rect 11698 9432 11704 9444
rect 10468 9404 11704 9432
rect 10468 9392 10474 9404
rect 11698 9392 11704 9404
rect 11756 9432 11762 9444
rect 11900 9432 11928 9463
rect 12158 9460 12164 9472
rect 12216 9500 12222 9512
rect 13372 9500 13400 9540
rect 12216 9472 13400 9500
rect 13909 9503 13967 9509
rect 12216 9460 12222 9472
rect 13909 9469 13921 9503
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 11756 9404 11928 9432
rect 11756 9392 11762 9404
rect 10134 9364 10140 9376
rect 7892 9336 10140 9364
rect 7892 9324 7898 9336
rect 10134 9324 10140 9336
rect 10192 9364 10198 9376
rect 11790 9364 11796 9376
rect 10192 9336 11796 9364
rect 10192 9324 10198 9336
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 11900 9364 11928 9404
rect 13170 9392 13176 9444
rect 13228 9432 13234 9444
rect 13924 9432 13952 9463
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 14274 9500 14280 9512
rect 14056 9472 14280 9500
rect 14056 9460 14062 9472
rect 14274 9460 14280 9472
rect 14332 9500 14338 9512
rect 15105 9503 15163 9509
rect 15105 9500 15117 9503
rect 14332 9472 15117 9500
rect 14332 9460 14338 9472
rect 15105 9469 15117 9472
rect 15151 9469 15163 9503
rect 15105 9463 15163 9469
rect 13228 9404 13952 9432
rect 13228 9392 13234 9404
rect 14016 9364 14044 9460
rect 15212 9432 15240 9540
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 16482 9568 16488 9580
rect 15841 9531 15899 9537
rect 15948 9540 16488 9568
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 15948 9500 15976 9540
rect 16482 9528 16488 9540
rect 16540 9528 16546 9580
rect 17880 9568 17908 9608
rect 18601 9605 18613 9639
rect 18647 9636 18659 9639
rect 21266 9636 21272 9648
rect 18647 9608 21272 9636
rect 18647 9605 18659 9608
rect 18601 9599 18659 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 21453 9639 21511 9645
rect 21453 9605 21465 9639
rect 21499 9636 21511 9639
rect 22370 9636 22376 9648
rect 21499 9608 22376 9636
rect 21499 9605 21511 9608
rect 21453 9599 21511 9605
rect 22370 9596 22376 9608
rect 22428 9596 22434 9648
rect 22738 9636 22744 9648
rect 22699 9608 22744 9636
rect 22738 9596 22744 9608
rect 22796 9596 22802 9648
rect 17696 9540 17908 9568
rect 16114 9500 16120 9512
rect 15436 9472 15976 9500
rect 16075 9472 16120 9500
rect 15436 9460 15442 9472
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 16390 9432 16396 9444
rect 15212 9404 16396 9432
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 16850 9392 16856 9444
rect 16908 9432 16914 9444
rect 16960 9432 16988 9463
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 17696 9500 17724 9540
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 19208 9540 19625 9568
rect 19208 9528 19214 9540
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 21818 9568 21824 9580
rect 19613 9531 19671 9537
rect 19904 9540 21824 9568
rect 19904 9512 19932 9540
rect 21818 9528 21824 9540
rect 21876 9528 21882 9580
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21968 9540 22017 9568
rect 21968 9528 21974 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9568 22707 9571
rect 23106 9568 23112 9580
rect 22695 9540 23112 9568
rect 22695 9537 22707 9540
rect 22649 9531 22707 9537
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9568 23351 9571
rect 24026 9568 24032 9580
rect 23339 9540 24032 9568
rect 23339 9537 23351 9540
rect 23293 9531 23351 9537
rect 24026 9528 24032 9540
rect 24084 9528 24090 9580
rect 24486 9568 24492 9580
rect 24447 9540 24492 9568
rect 24486 9528 24492 9540
rect 24544 9528 24550 9580
rect 24578 9528 24584 9580
rect 24636 9568 24642 9580
rect 25777 9571 25835 9577
rect 25777 9568 25789 9571
rect 24636 9540 25789 9568
rect 24636 9528 24642 9540
rect 25777 9537 25789 9540
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 17460 9472 17724 9500
rect 17460 9460 17466 9472
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18104 9472 18521 9500
rect 18104 9460 18110 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 18785 9503 18843 9509
rect 18785 9469 18797 9503
rect 18831 9469 18843 9503
rect 19886 9500 19892 9512
rect 19799 9472 19892 9500
rect 18785 9463 18843 9469
rect 16908 9404 16988 9432
rect 16908 9392 16914 9404
rect 17770 9392 17776 9444
rect 17828 9432 17834 9444
rect 18800 9432 18828 9463
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 20530 9460 20536 9512
rect 20588 9500 20594 9512
rect 20809 9503 20867 9509
rect 20809 9500 20821 9503
rect 20588 9472 20821 9500
rect 20588 9460 20594 9472
rect 20809 9469 20821 9472
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 20993 9503 21051 9509
rect 20993 9469 21005 9503
rect 21039 9500 21051 9503
rect 23385 9503 23443 9509
rect 23385 9500 23397 9503
rect 21039 9472 23397 9500
rect 21039 9469 21051 9472
rect 20993 9463 21051 9469
rect 23385 9469 23397 9472
rect 23431 9469 23443 9503
rect 23385 9463 23443 9469
rect 24673 9503 24731 9509
rect 24673 9469 24685 9503
rect 24719 9469 24731 9503
rect 24673 9463 24731 9469
rect 17828 9404 18828 9432
rect 17828 9392 17834 9404
rect 18874 9392 18880 9444
rect 18932 9432 18938 9444
rect 23198 9432 23204 9444
rect 18932 9404 23204 9432
rect 18932 9392 18938 9404
rect 23198 9392 23204 9404
rect 23256 9392 23262 9444
rect 24688 9432 24716 9463
rect 25593 9435 25651 9441
rect 25593 9432 25605 9435
rect 24688 9404 25605 9432
rect 25593 9401 25605 9404
rect 25639 9401 25651 9435
rect 25593 9395 25651 9401
rect 11900 9336 14044 9364
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 15746 9364 15752 9376
rect 14516 9336 15752 9364
rect 14516 9324 14522 9336
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 15930 9324 15936 9376
rect 15988 9364 15994 9376
rect 19886 9364 19892 9376
rect 15988 9336 19892 9364
rect 15988 9324 15994 9336
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 22094 9364 22100 9376
rect 22055 9336 22100 9364
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 24854 9364 24860 9376
rect 24815 9336 24860 9364
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2590 9160 2596 9172
rect 2551 9132 2596 9160
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 5629 9163 5687 9169
rect 2740 9132 4752 9160
rect 2740 9120 2746 9132
rect 2130 9052 2136 9104
rect 2188 9092 2194 9104
rect 3329 9095 3387 9101
rect 3329 9092 3341 9095
rect 2188 9064 3341 9092
rect 2188 9052 2194 9064
rect 3329 9061 3341 9064
rect 3375 9061 3387 9095
rect 3329 9055 3387 9061
rect 3602 9052 3608 9104
rect 3660 9092 3666 9104
rect 4614 9092 4620 9104
rect 3660 9064 4620 9092
rect 3660 9052 3666 9064
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 4724 9092 4752 9132
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 7742 9160 7748 9172
rect 5675 9132 7748 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 9401 9163 9459 9169
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 11514 9160 11520 9172
rect 9447 9132 11520 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 12176 9132 12357 9160
rect 5902 9092 5908 9104
rect 4724 9064 5908 9092
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 7929 9095 7987 9101
rect 7929 9092 7941 9095
rect 7616 9064 7941 9092
rect 7616 9052 7622 9064
rect 7929 9061 7941 9064
rect 7975 9061 7987 9095
rect 12176 9092 12204 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 16040 9132 18644 9160
rect 7929 9055 7987 9061
rect 11992 9064 12204 9092
rect 4706 9024 4712 9036
rect 2516 8996 3188 9024
rect 4667 8996 4712 9024
rect 2516 8968 2544 8996
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1544 8928 1593 8956
rect 1544 8916 1550 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 2498 8916 2504 8968
rect 2556 8916 2562 8968
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 2832 8928 2877 8956
rect 2832 8916 2838 8928
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 3160 8820 3188 8996
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 6454 9024 6460 9036
rect 6415 8996 6460 9024
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 6604 8996 10272 9024
rect 6604 8984 6610 8996
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 4890 8956 4896 8968
rect 3283 8928 4896 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 3973 8891 4031 8897
rect 3973 8857 3985 8891
rect 4019 8888 4031 8891
rect 4614 8888 4620 8900
rect 4019 8860 4620 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 5552 8888 5580 8919
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 6181 8959 6239 8965
rect 6181 8956 6193 8959
rect 5960 8928 6193 8956
rect 5960 8916 5966 8928
rect 6181 8925 6193 8928
rect 6227 8925 6239 8959
rect 8018 8956 8024 8968
rect 7590 8928 8024 8956
rect 6181 8919 6239 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8956 9367 8959
rect 9858 8956 9864 8968
rect 9355 8928 9864 8956
rect 9355 8925 9367 8928
rect 9309 8919 9367 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 5626 8888 5632 8900
rect 5539 8860 5632 8888
rect 5626 8848 5632 8860
rect 5684 8888 5690 8900
rect 6730 8888 6736 8900
rect 5684 8860 6736 8888
rect 5684 8848 5690 8860
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 7742 8848 7748 8900
rect 7800 8888 7806 8900
rect 10244 8888 10272 8996
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 10468 8996 10609 9024
rect 10468 8984 10474 8996
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 10962 9024 10968 9036
rect 10919 8996 10968 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 11992 9024 12020 9064
rect 14274 9024 14280 9036
rect 11664 8996 12020 9024
rect 14235 8996 14280 9024
rect 11664 8984 11670 8996
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 14918 8984 14924 9036
rect 14976 9024 14982 9036
rect 16040 9033 16068 9132
rect 16482 9052 16488 9104
rect 16540 9092 16546 9104
rect 18506 9092 18512 9104
rect 16540 9064 18512 9092
rect 16540 9052 16546 9064
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 18616 9092 18644 9132
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 18966 9160 18972 9172
rect 18748 9132 18972 9160
rect 18748 9120 18754 9132
rect 18966 9120 18972 9132
rect 19024 9160 19030 9172
rect 19978 9160 19984 9172
rect 19024 9132 19984 9160
rect 19024 9120 19030 9132
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 20714 9160 20720 9172
rect 20675 9132 20720 9160
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 23842 9160 23848 9172
rect 23803 9132 23848 9160
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 24578 9160 24584 9172
rect 24539 9132 24584 9160
rect 24578 9120 24584 9132
rect 24636 9120 24642 9172
rect 25498 9120 25504 9172
rect 25556 9160 25562 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 25556 9132 29837 9160
rect 25556 9120 25562 9132
rect 29825 9129 29837 9132
rect 29871 9129 29883 9163
rect 29825 9123 29883 9129
rect 18874 9092 18880 9104
rect 18616 9064 18880 9092
rect 18874 9052 18880 9064
rect 18932 9052 18938 9104
rect 22646 9092 22652 9104
rect 19628 9064 22652 9092
rect 19521 9039 19579 9045
rect 16025 9027 16083 9033
rect 16025 9024 16037 9027
rect 14976 8996 16037 9024
rect 14976 8984 14982 8996
rect 16025 8993 16037 8996
rect 16071 8993 16083 9027
rect 16025 8987 16083 8993
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 9024 17095 9027
rect 18782 9024 18788 9036
rect 17083 8996 18788 9024
rect 17083 8993 17095 8996
rect 17037 8987 17095 8993
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 19521 9005 19533 9039
rect 19567 9036 19579 9039
rect 19628 9036 19656 9064
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 19567 9008 19656 9036
rect 19978 9024 19984 9036
rect 19567 9005 19579 9008
rect 19521 8999 19579 9005
rect 19939 8996 19984 9024
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 22557 9027 22615 9033
rect 22557 9024 22569 9027
rect 20956 8996 22569 9024
rect 20956 8984 20962 8996
rect 22557 8993 22569 8996
rect 22603 8993 22615 9027
rect 22557 8987 22615 8993
rect 23382 8984 23388 9036
rect 23440 9024 23446 9036
rect 23440 8996 24808 9024
rect 23440 8984 23446 8996
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 13262 8956 13268 8968
rect 12400 8928 13268 8956
rect 12400 8916 12406 8928
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13722 8956 13728 8968
rect 13464 8928 13728 8956
rect 13464 8888 13492 8928
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 13998 8916 14004 8968
rect 14056 8916 14062 8968
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16264 8928 16865 8956
rect 16264 8916 16270 8928
rect 16853 8925 16865 8928
rect 16899 8956 16911 8959
rect 17770 8956 17776 8968
rect 16899 8928 17776 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 18690 8916 18696 8968
rect 18748 8956 18754 8968
rect 18748 8928 18793 8956
rect 18748 8916 18754 8928
rect 20346 8916 20352 8968
rect 20404 8956 20410 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20404 8928 20637 8956
rect 20404 8916 20410 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 22465 8959 22523 8965
rect 22465 8925 22477 8959
rect 22511 8925 22523 8959
rect 22465 8919 22523 8925
rect 7800 8860 10088 8888
rect 10244 8860 11362 8888
rect 12360 8860 13492 8888
rect 13541 8891 13599 8897
rect 7800 8848 7806 8860
rect 8754 8820 8760 8832
rect 3160 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9950 8820 9956 8832
rect 9911 8792 9956 8820
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10060 8820 10088 8860
rect 12360 8820 12388 8860
rect 13541 8857 13553 8891
rect 13587 8888 13599 8891
rect 14016 8888 14044 8916
rect 14550 8888 14556 8900
rect 13587 8860 14044 8888
rect 14511 8860 14556 8888
rect 13587 8857 13599 8860
rect 13541 8851 13599 8857
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 15194 8848 15200 8900
rect 15252 8848 15258 8900
rect 16574 8888 16580 8900
rect 15856 8860 16580 8888
rect 10060 8792 12388 8820
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 15856 8820 15884 8860
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 18046 8888 18052 8900
rect 16776 8860 18052 8888
rect 12584 8792 15884 8820
rect 12584 8780 12590 8792
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 16776 8820 16804 8860
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 18138 8848 18144 8900
rect 18196 8888 18202 8900
rect 19613 8891 19671 8897
rect 18196 8860 18241 8888
rect 18616 8860 19564 8888
rect 18196 8848 18202 8860
rect 17494 8820 17500 8832
rect 15988 8792 16804 8820
rect 17455 8792 17500 8820
rect 15988 8780 15994 8792
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 18616 8820 18644 8860
rect 17644 8792 18644 8820
rect 17644 8780 17650 8792
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 19334 8820 19340 8832
rect 18932 8792 19340 8820
rect 18932 8780 18938 8792
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19536 8820 19564 8860
rect 19613 8857 19625 8891
rect 19659 8888 19671 8891
rect 20806 8888 20812 8900
rect 19659 8860 20812 8888
rect 19659 8857 19671 8860
rect 19613 8851 19671 8857
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 21361 8891 21419 8897
rect 21361 8888 21373 8891
rect 21232 8860 21373 8888
rect 21232 8848 21238 8860
rect 21361 8857 21373 8860
rect 21407 8857 21419 8891
rect 21361 8851 21419 8857
rect 21450 8848 21456 8900
rect 21508 8888 21514 8900
rect 21508 8860 21553 8888
rect 21508 8848 21514 8860
rect 21726 8848 21732 8900
rect 21784 8888 21790 8900
rect 22005 8891 22063 8897
rect 22005 8888 22017 8891
rect 21784 8860 22017 8888
rect 21784 8848 21790 8860
rect 22005 8857 22017 8860
rect 22051 8857 22063 8891
rect 22005 8851 22063 8857
rect 21910 8820 21916 8832
rect 19536 8792 21916 8820
rect 21910 8780 21916 8792
rect 21968 8820 21974 8832
rect 22480 8820 22508 8919
rect 22738 8916 22744 8968
rect 22796 8956 22802 8968
rect 23109 8959 23167 8965
rect 23109 8956 23121 8959
rect 22796 8928 23121 8956
rect 22796 8916 22802 8928
rect 23109 8925 23121 8928
rect 23155 8925 23167 8959
rect 23109 8919 23167 8925
rect 23753 8959 23811 8965
rect 23753 8925 23765 8959
rect 23799 8956 23811 8959
rect 23934 8956 23940 8968
rect 23799 8928 23940 8956
rect 23799 8925 23811 8928
rect 23753 8919 23811 8925
rect 23934 8916 23940 8928
rect 23992 8916 23998 8968
rect 24780 8965 24808 8996
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8925 24823 8959
rect 25222 8956 25228 8968
rect 25183 8928 25228 8956
rect 24765 8919 24823 8925
rect 25222 8916 25228 8928
rect 25280 8916 25286 8968
rect 29733 8959 29791 8965
rect 29733 8925 29745 8959
rect 29779 8956 29791 8959
rect 30742 8956 30748 8968
rect 29779 8928 30748 8956
rect 29779 8925 29791 8928
rect 29733 8919 29791 8925
rect 30742 8916 30748 8928
rect 30800 8916 30806 8968
rect 21968 8792 22508 8820
rect 21968 8780 21974 8792
rect 22554 8780 22560 8832
rect 22612 8820 22618 8832
rect 23201 8823 23259 8829
rect 23201 8820 23213 8823
rect 22612 8792 23213 8820
rect 22612 8780 22618 8792
rect 23201 8789 23213 8792
rect 23247 8789 23259 8823
rect 25314 8820 25320 8832
rect 25275 8792 25320 8820
rect 23201 8783 23259 8789
rect 25314 8780 25320 8792
rect 25372 8780 25378 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1765 8619 1823 8625
rect 1765 8616 1777 8619
rect 1452 8588 1777 8616
rect 1452 8576 1458 8588
rect 1765 8585 1777 8588
rect 1811 8585 1823 8619
rect 2866 8616 2872 8628
rect 1765 8579 1823 8585
rect 1964 8588 2872 8616
rect 1964 8489 1992 8588
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 5261 8619 5319 8625
rect 5261 8585 5273 8619
rect 5307 8616 5319 8619
rect 7742 8616 7748 8628
rect 5307 8588 7748 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 9398 8616 9404 8628
rect 8036 8588 9404 8616
rect 2685 8551 2743 8557
rect 2685 8517 2697 8551
rect 2731 8548 2743 8551
rect 2958 8548 2964 8560
rect 2731 8520 2964 8548
rect 2731 8517 2743 8520
rect 2685 8511 2743 8517
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 4706 8548 4712 8560
rect 3910 8520 4712 8548
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 6641 8551 6699 8557
rect 5592 8520 6592 8548
rect 5592 8508 5598 8520
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 6564 8489 6592 8520
rect 6641 8517 6653 8551
rect 6687 8548 6699 8551
rect 8036 8548 8064 8588
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 13262 8616 13268 8628
rect 10008 8588 13268 8616
rect 10008 8576 10014 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 13964 8588 16221 8616
rect 13964 8576 13970 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 17494 8616 17500 8628
rect 17455 8588 17500 8616
rect 16209 8579 16267 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 19702 8616 19708 8628
rect 17920 8588 19708 8616
rect 17920 8576 17926 8588
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20990 8616 20996 8628
rect 19812 8588 20996 8616
rect 6687 8520 8064 8548
rect 6687 8517 6699 8520
rect 6641 8511 6699 8517
rect 8478 8508 8484 8560
rect 8536 8508 8542 8560
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 10137 8551 10195 8557
rect 10137 8548 10149 8551
rect 9272 8520 10149 8548
rect 9272 8508 9278 8520
rect 10137 8517 10149 8520
rect 10183 8517 10195 8551
rect 12342 8548 12348 8560
rect 10137 8511 10195 8517
rect 10704 8520 12348 8548
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 4028 8452 5181 8480
rect 4028 8440 4034 8452
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5169 8443 5227 8449
rect 5644 8452 5825 8480
rect 2222 8372 2228 8424
rect 2280 8412 2286 8424
rect 2409 8415 2467 8421
rect 2409 8412 2421 8415
rect 2280 8384 2421 8412
rect 2280 8372 2286 8384
rect 2409 8381 2421 8384
rect 2455 8381 2467 8415
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 2409 8375 2467 8381
rect 2516 8384 4169 8412
rect 1302 8304 1308 8356
rect 1360 8344 1366 8356
rect 2516 8344 2544 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4982 8372 4988 8424
rect 5040 8412 5046 8424
rect 5534 8412 5540 8424
rect 5040 8384 5540 8412
rect 5040 8372 5046 8384
rect 5534 8372 5540 8384
rect 5592 8412 5598 8424
rect 5644 8412 5672 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 10045 8483 10103 8489
rect 6549 8443 6607 8449
rect 9232 8452 9996 8480
rect 5592 8384 5672 8412
rect 5592 8372 5598 8384
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 5776 8384 5917 8412
rect 5776 8372 5782 8384
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 7466 8412 7472 8424
rect 7379 8384 7472 8412
rect 5905 8375 5963 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 9232 8412 9260 8452
rect 7791 8384 9260 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9364 8384 9505 8412
rect 9364 8372 9370 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9968 8412 9996 8452
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10410 8480 10416 8492
rect 10091 8452 10416 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10704 8489 10732 8520
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 12986 8508 12992 8560
rect 13044 8508 13050 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 14645 8551 14703 8557
rect 14645 8548 14657 8551
rect 13596 8520 14657 8548
rect 13596 8508 13602 8520
rect 14645 8517 14657 8520
rect 14691 8517 14703 8551
rect 14645 8511 14703 8517
rect 14734 8508 14740 8560
rect 14792 8548 14798 8560
rect 14792 8520 14837 8548
rect 14792 8508 14798 8520
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 15160 8520 16160 8548
rect 15160 8508 15166 8520
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 10965 8483 11023 8489
rect 10965 8480 10977 8483
rect 10836 8452 10977 8480
rect 10836 8440 10842 8452
rect 10965 8449 10977 8452
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11698 8480 11704 8492
rect 11204 8452 11704 8480
rect 11204 8440 11210 8452
rect 11698 8440 11704 8452
rect 11756 8480 11762 8492
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11756 8452 11989 8480
rect 11756 8440 11762 8452
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 14458 8480 14464 8492
rect 11977 8443 12035 8449
rect 14016 8452 14464 8480
rect 10870 8412 10876 8424
rect 9968 8384 10876 8412
rect 9493 8375 9551 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 11296 8384 12265 8412
rect 11296 8372 11302 8384
rect 12253 8381 12265 8384
rect 12299 8381 12311 8415
rect 12253 8375 12311 8381
rect 12710 8372 12716 8424
rect 12768 8412 12774 8424
rect 14016 8421 14044 8452
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 16132 8489 16160 8520
rect 18046 8508 18052 8560
rect 18104 8548 18110 8560
rect 18141 8551 18199 8557
rect 18141 8548 18153 8551
rect 18104 8520 18153 8548
rect 18104 8508 18110 8520
rect 18141 8517 18153 8520
rect 18187 8517 18199 8551
rect 18141 8511 18199 8517
rect 18598 8508 18604 8560
rect 18656 8548 18662 8560
rect 18656 8520 19334 8548
rect 18656 8508 18662 8520
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16816 8452 16865 8480
rect 16816 8440 16822 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 17586 8480 17592 8492
rect 16853 8443 16911 8449
rect 16960 8452 17592 8480
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 12768 8384 14013 8412
rect 12768 8372 12774 8384
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 15102 8412 15108 8424
rect 14148 8384 15108 8412
rect 14148 8372 14154 8384
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 15657 8415 15715 8421
rect 15657 8412 15669 8415
rect 15620 8384 15669 8412
rect 15620 8372 15626 8384
rect 15657 8381 15669 8384
rect 15703 8412 15715 8415
rect 15746 8412 15752 8424
rect 15703 8384 15752 8412
rect 15703 8381 15715 8384
rect 15657 8375 15715 8381
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 1360 8316 2544 8344
rect 1360 8304 1366 8316
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 7374 8344 7380 8356
rect 3752 8316 7380 8344
rect 3752 8304 3758 8316
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 6546 8276 6552 8288
rect 5776 8248 6552 8276
rect 5776 8236 5782 8248
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 7484 8276 7512 8372
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 10502 8344 10508 8356
rect 9180 8316 10508 8344
rect 9180 8304 9186 8316
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 16960 8344 16988 8452
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 19306 8480 19334 8520
rect 19812 8480 19840 8588
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 22094 8616 22100 8628
rect 21100 8588 22100 8616
rect 20073 8551 20131 8557
rect 20073 8517 20085 8551
rect 20119 8548 20131 8551
rect 21100 8548 21128 8588
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 25133 8619 25191 8625
rect 25133 8616 25145 8619
rect 22848 8588 25145 8616
rect 21358 8548 21364 8560
rect 20119 8520 21128 8548
rect 21319 8520 21364 8548
rect 20119 8517 20131 8520
rect 20073 8511 20131 8517
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 21450 8508 21456 8560
rect 21508 8548 21514 8560
rect 22848 8548 22876 8588
rect 25133 8585 25145 8588
rect 25179 8585 25191 8619
rect 25133 8579 25191 8585
rect 33042 8576 33048 8628
rect 33100 8616 33106 8628
rect 38105 8619 38163 8625
rect 38105 8616 38117 8619
rect 33100 8588 38117 8616
rect 33100 8576 33106 8588
rect 38105 8585 38117 8588
rect 38151 8585 38163 8619
rect 38105 8579 38163 8585
rect 21508 8520 22876 8548
rect 22940 8520 31754 8548
rect 21508 8508 21514 8520
rect 19306 8452 19840 8480
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20714 8480 20720 8492
rect 20671 8452 20720 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 21082 8440 21088 8492
rect 21140 8480 21146 8492
rect 21177 8483 21235 8489
rect 21177 8480 21189 8483
rect 21140 8452 21189 8480
rect 21140 8440 21146 8452
rect 21177 8449 21189 8452
rect 21223 8449 21235 8483
rect 22002 8480 22008 8492
rect 21963 8452 22008 8480
rect 21177 8443 21235 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 17037 8415 17095 8421
rect 17037 8381 17049 8415
rect 17083 8381 17095 8415
rect 17037 8375 17095 8381
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18230 8412 18236 8424
rect 18095 8384 18236 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 13780 8316 16988 8344
rect 17052 8344 17080 8375
rect 18230 8372 18236 8384
rect 18288 8412 18294 8424
rect 18506 8412 18512 8424
rect 18288 8384 18512 8412
rect 18288 8372 18294 8384
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 18598 8372 18604 8424
rect 18656 8412 18662 8424
rect 18656 8384 18701 8412
rect 18656 8372 18662 8384
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 19794 8412 19800 8424
rect 19116 8384 19800 8412
rect 19116 8372 19122 8384
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20346 8412 20352 8424
rect 20027 8384 20352 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 20898 8412 20904 8424
rect 20456 8384 20904 8412
rect 20456 8344 20484 8384
rect 20898 8372 20904 8384
rect 20956 8372 20962 8424
rect 20990 8372 20996 8424
rect 21048 8412 21054 8424
rect 22940 8412 22968 8520
rect 23382 8440 23388 8492
rect 23440 8480 23446 8492
rect 24121 8483 24179 8489
rect 24121 8480 24133 8483
rect 23440 8452 24133 8480
rect 23440 8440 23446 8452
rect 24121 8449 24133 8452
rect 24167 8449 24179 8483
rect 25038 8480 25044 8492
rect 24999 8452 25044 8480
rect 24121 8443 24179 8449
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 31726 8480 31754 8520
rect 32953 8483 33011 8489
rect 32953 8480 32965 8483
rect 31726 8452 32965 8480
rect 25685 8443 25743 8449
rect 32953 8449 32965 8452
rect 32999 8449 33011 8483
rect 38286 8480 38292 8492
rect 38247 8452 38292 8480
rect 32953 8443 33011 8449
rect 21048 8384 22968 8412
rect 23017 8415 23075 8421
rect 21048 8372 21054 8384
rect 23017 8381 23029 8415
rect 23063 8381 23075 8415
rect 23017 8375 23075 8381
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8412 23259 8415
rect 24213 8415 24271 8421
rect 24213 8412 24225 8415
rect 23247 8384 24225 8412
rect 23247 8381 23259 8384
rect 23201 8375 23259 8381
rect 24213 8381 24225 8384
rect 24259 8381 24271 8415
rect 24213 8375 24271 8381
rect 17052 8316 20484 8344
rect 13780 8304 13786 8316
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 22097 8347 22155 8353
rect 22097 8344 22109 8347
rect 20588 8316 22109 8344
rect 20588 8304 20594 8316
rect 22097 8313 22109 8316
rect 22143 8313 22155 8347
rect 22097 8307 22155 8313
rect 22370 8304 22376 8356
rect 22428 8344 22434 8356
rect 23032 8344 23060 8375
rect 22428 8316 23060 8344
rect 23661 8347 23719 8353
rect 22428 8304 22434 8316
rect 23661 8313 23673 8347
rect 23707 8344 23719 8347
rect 24854 8344 24860 8356
rect 23707 8316 24860 8344
rect 23707 8313 23719 8316
rect 23661 8307 23719 8313
rect 24854 8304 24860 8316
rect 24912 8344 24918 8356
rect 25700 8344 25728 8443
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 24912 8316 25728 8344
rect 25777 8347 25835 8353
rect 24912 8304 24918 8316
rect 25777 8313 25789 8347
rect 25823 8344 25835 8347
rect 26142 8344 26148 8356
rect 25823 8316 26148 8344
rect 25823 8313 25835 8316
rect 25777 8307 25835 8313
rect 26142 8304 26148 8316
rect 26200 8304 26206 8356
rect 33045 8347 33103 8353
rect 33045 8313 33057 8347
rect 33091 8344 33103 8347
rect 34422 8344 34428 8356
rect 33091 8316 34428 8344
rect 33091 8313 33103 8316
rect 33045 8307 33103 8313
rect 34422 8304 34428 8316
rect 34480 8304 34486 8356
rect 9140 8276 9168 8304
rect 7484 8248 9168 8276
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 10226 8276 10232 8288
rect 9364 8248 10232 8276
rect 9364 8236 9370 8248
rect 10226 8236 10232 8248
rect 10284 8276 10290 8288
rect 10410 8276 10416 8288
rect 10284 8248 10416 8276
rect 10284 8236 10290 8248
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 15194 8276 15200 8288
rect 11296 8248 15200 8276
rect 11296 8236 11302 8248
rect 15194 8236 15200 8248
rect 15252 8236 15258 8288
rect 16482 8236 16488 8288
rect 16540 8276 16546 8288
rect 24762 8276 24768 8288
rect 16540 8248 24768 8276
rect 16540 8236 16546 8248
rect 24762 8236 24768 8248
rect 24820 8236 24826 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 1728 8044 2973 8072
rect 1728 8032 1734 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 13538 8072 13544 8084
rect 2961 8035 3019 8041
rect 5736 8044 13544 8072
rect 4522 7964 4528 8016
rect 4580 8004 4586 8016
rect 5626 8004 5632 8016
rect 4580 7976 5632 8004
rect 4580 7964 4586 7976
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 934 7896 940 7948
rect 992 7936 998 7948
rect 1857 7939 1915 7945
rect 1857 7936 1869 7939
rect 992 7908 1869 7936
rect 992 7896 998 7908
rect 1857 7905 1869 7908
rect 1903 7905 1915 7939
rect 1857 7899 1915 7905
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 4982 7936 4988 7948
rect 3844 7908 4988 7936
rect 3844 7896 3850 7908
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 2866 7868 2872 7880
rect 2827 7840 2872 7868
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4632 7877 4660 7908
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5736 7936 5764 8044
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14240 8044 16068 8072
rect 14240 8032 14246 8044
rect 16040 8016 16068 8044
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 18046 8072 18052 8084
rect 16448 8044 18052 8072
rect 16448 8032 16454 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18230 8032 18236 8084
rect 18288 8072 18294 8084
rect 18288 8044 20208 8072
rect 18288 8032 18294 8044
rect 7650 8004 7656 8016
rect 7611 7976 7656 8004
rect 7650 7964 7656 7976
rect 7708 7964 7714 8016
rect 10873 8007 10931 8013
rect 8128 7976 9260 8004
rect 5123 7908 5764 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 8128 7936 8156 7976
rect 6696 7908 8156 7936
rect 6696 7896 6702 7908
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8846 7936 8852 7948
rect 8352 7908 8852 7936
rect 8352 7896 8358 7908
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 9122 7936 9128 7948
rect 9083 7908 9128 7936
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 9232 7936 9260 7976
rect 10873 7973 10885 8007
rect 10919 8004 10931 8007
rect 10962 8004 10968 8016
rect 10919 7976 10968 8004
rect 10919 7973 10931 7976
rect 10873 7967 10931 7973
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 16022 8004 16028 8016
rect 15935 7976 16028 8004
rect 16022 7964 16028 7976
rect 16080 8004 16086 8016
rect 16080 7976 17908 8004
rect 16080 7964 16086 7976
rect 11146 7936 11152 7948
rect 9232 7908 11152 7936
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 11609 7939 11667 7945
rect 11609 7905 11621 7939
rect 11655 7936 11667 7939
rect 11698 7936 11704 7948
rect 11655 7908 11704 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7936 13415 7939
rect 13630 7936 13636 7948
rect 13403 7908 13636 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 15194 7936 15200 7948
rect 15155 7908 15200 7936
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7936 16727 7939
rect 17494 7936 17500 7948
rect 16715 7908 17500 7936
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 17770 7936 17776 7948
rect 17644 7908 17776 7936
rect 17644 7896 17650 7908
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 17880 7936 17908 7976
rect 18414 7964 18420 8016
rect 18472 7964 18478 8016
rect 19705 8007 19763 8013
rect 19705 7973 19717 8007
rect 19751 8004 19763 8007
rect 20070 8004 20076 8016
rect 19751 7976 20076 8004
rect 19751 7973 19763 7976
rect 19705 7967 19763 7973
rect 20070 7964 20076 7976
rect 20128 7964 20134 8016
rect 20180 8004 20208 8044
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 20714 8072 20720 8084
rect 20312 8044 20720 8072
rect 20312 8032 20318 8044
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 23385 8075 23443 8081
rect 23385 8072 23397 8075
rect 20864 8044 23397 8072
rect 20864 8032 20870 8044
rect 23385 8041 23397 8044
rect 23431 8041 23443 8075
rect 31386 8072 31392 8084
rect 31347 8044 31392 8072
rect 23385 8035 23443 8041
rect 31386 8032 31392 8044
rect 31444 8032 31450 8084
rect 24673 8007 24731 8013
rect 24673 8004 24685 8007
rect 20180 7976 24685 8004
rect 24673 7973 24685 7976
rect 24719 7973 24731 8007
rect 38105 8007 38163 8013
rect 38105 8004 38117 8007
rect 24673 7967 24731 7973
rect 31726 7976 38117 8004
rect 18432 7936 18460 7964
rect 17880 7908 18460 7936
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7868 4767 7871
rect 5718 7868 5724 7880
rect 4755 7840 5724 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 6181 7803 6239 7809
rect 6181 7769 6193 7803
rect 6227 7800 6239 7803
rect 6454 7800 6460 7812
rect 6227 7772 6460 7800
rect 6227 7769 6239 7772
rect 6181 7763 6239 7769
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 8202 7800 8208 7812
rect 7406 7772 8208 7800
rect 4065 7735 4123 7741
rect 4065 7701 4077 7735
rect 4111 7732 4123 7735
rect 4982 7732 4988 7744
rect 4111 7704 4988 7732
rect 4111 7701 4123 7704
rect 4065 7695 4123 7701
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 7484 7732 7512 7772
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 8404 7800 8432 7831
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11112 7840 11345 7868
rect 11112 7828 11118 7840
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7868 15899 7871
rect 16482 7868 16488 7880
rect 15887 7840 16488 7868
rect 15887 7837 15899 7840
rect 15841 7831 15899 7837
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 18156 7877 18184 7908
rect 19794 7896 19800 7948
rect 19852 7936 19858 7948
rect 20346 7936 20352 7948
rect 19852 7908 20208 7936
rect 20259 7908 20352 7936
rect 19852 7896 19858 7908
rect 20180 7880 20208 7908
rect 20346 7896 20352 7908
rect 20404 7936 20410 7948
rect 20714 7936 20720 7948
rect 20404 7908 20720 7936
rect 20404 7896 20410 7908
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 20806 7896 20812 7948
rect 20864 7936 20870 7948
rect 20864 7908 20909 7936
rect 20864 7896 20870 7908
rect 21174 7896 21180 7948
rect 21232 7936 21238 7948
rect 21545 7939 21603 7945
rect 21545 7936 21557 7939
rect 21232 7908 21557 7936
rect 21232 7896 21238 7908
rect 21545 7905 21557 7908
rect 21591 7905 21603 7939
rect 21545 7899 21603 7905
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 24026 7936 24032 7948
rect 21876 7908 24032 7936
rect 21876 7896 21882 7908
rect 24026 7896 24032 7908
rect 24084 7896 24090 7948
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18322 7828 18328 7880
rect 18380 7868 18386 7880
rect 18417 7871 18475 7877
rect 18417 7868 18429 7871
rect 18380 7840 18429 7868
rect 18380 7828 18386 7840
rect 18417 7837 18429 7840
rect 18463 7868 18475 7871
rect 20070 7868 20076 7880
rect 18463 7840 20076 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 20162 7828 20168 7880
rect 20220 7828 20226 7880
rect 22646 7868 22652 7880
rect 22607 7840 22652 7868
rect 22646 7828 22652 7840
rect 22704 7828 22710 7880
rect 23198 7828 23204 7880
rect 23256 7868 23262 7880
rect 23293 7871 23351 7877
rect 23293 7868 23305 7871
rect 23256 7840 23305 7868
rect 23256 7828 23262 7840
rect 23293 7837 23305 7840
rect 23339 7837 23351 7871
rect 23293 7831 23351 7837
rect 23382 7828 23388 7880
rect 23440 7868 23446 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 23440 7840 24593 7868
rect 23440 7828 23446 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 31297 7871 31355 7877
rect 31297 7837 31309 7871
rect 31343 7868 31355 7871
rect 31726 7868 31754 7976
rect 38105 7973 38117 7976
rect 38151 7973 38163 8007
rect 38105 7967 38163 7973
rect 31343 7840 31754 7868
rect 31343 7837 31355 7840
rect 31297 7831 31355 7837
rect 34422 7828 34428 7880
rect 34480 7868 34486 7880
rect 35713 7871 35771 7877
rect 35713 7868 35725 7871
rect 34480 7840 35725 7868
rect 34480 7828 34486 7840
rect 35713 7837 35725 7840
rect 35759 7837 35771 7871
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 35713 7831 35771 7837
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 9306 7800 9312 7812
rect 8404 7772 9312 7800
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 9398 7760 9404 7812
rect 9456 7800 9462 7812
rect 10962 7800 10968 7812
rect 9456 7772 9501 7800
rect 10626 7772 10968 7800
rect 9456 7760 9462 7772
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 14737 7803 14795 7809
rect 11532 7772 12098 7800
rect 5675 7704 7512 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 8481 7735 8539 7741
rect 8481 7732 8493 7735
rect 8444 7704 8493 7732
rect 8444 7692 8450 7704
rect 8481 7701 8493 7704
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 11532 7732 11560 7772
rect 14737 7769 14749 7803
rect 14783 7769 14795 7803
rect 14737 7763 14795 7769
rect 14829 7803 14887 7809
rect 14829 7769 14841 7803
rect 14875 7800 14887 7803
rect 16761 7803 16819 7809
rect 14875 7772 16712 7800
rect 14875 7769 14887 7772
rect 14829 7763 14887 7769
rect 8720 7704 11560 7732
rect 8720 7692 8726 7704
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 14752 7732 14780 7763
rect 16574 7732 16580 7744
rect 14608 7704 16580 7732
rect 14608 7692 14614 7704
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 16684 7732 16712 7772
rect 16761 7769 16773 7803
rect 16807 7800 16819 7803
rect 17862 7800 17868 7812
rect 16807 7772 17868 7800
rect 16807 7769 16819 7772
rect 16761 7763 16819 7769
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 19521 7803 19579 7809
rect 19521 7769 19533 7803
rect 19567 7800 19579 7803
rect 20346 7800 20352 7812
rect 19567 7772 20352 7800
rect 19567 7769 19579 7772
rect 19521 7763 19579 7769
rect 20346 7760 20352 7772
rect 20404 7760 20410 7812
rect 20441 7803 20499 7809
rect 20441 7769 20453 7803
rect 20487 7769 20499 7803
rect 20441 7763 20499 7769
rect 17494 7732 17500 7744
rect 16684 7704 17500 7732
rect 17494 7692 17500 7704
rect 17552 7692 17558 7744
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 20162 7732 20168 7744
rect 18012 7704 20168 7732
rect 18012 7692 18018 7704
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 20456 7732 20484 7763
rect 21634 7760 21640 7812
rect 21692 7800 21698 7812
rect 21692 7772 21737 7800
rect 21692 7760 21698 7772
rect 21818 7760 21824 7812
rect 21876 7800 21882 7812
rect 22189 7803 22247 7809
rect 22189 7800 22201 7803
rect 21876 7772 22201 7800
rect 21876 7760 21882 7772
rect 22189 7769 22201 7772
rect 22235 7769 22247 7803
rect 22189 7763 22247 7769
rect 22554 7732 22560 7744
rect 20456 7704 22560 7732
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 35529 7735 35587 7741
rect 35529 7701 35541 7735
rect 35575 7732 35587 7735
rect 38010 7732 38016 7744
rect 35575 7704 38016 7732
rect 35575 7701 35587 7704
rect 35529 7695 35587 7701
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 4798 7528 4804 7540
rect 2746 7500 4804 7528
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7460 2559 7463
rect 2746 7460 2774 7500
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 8386 7528 8392 7540
rect 5868 7500 8392 7528
rect 5868 7488 5874 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 13170 7528 13176 7540
rect 9456 7500 13176 7528
rect 9456 7488 9462 7500
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 18322 7528 18328 7540
rect 14148 7500 18328 7528
rect 14148 7488 14154 7500
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 20898 7528 20904 7540
rect 19444 7500 20904 7528
rect 5368 7460 5396 7488
rect 2547 7432 2774 7460
rect 3726 7432 5396 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 7285 7463 7343 7469
rect 7285 7460 7297 7463
rect 5960 7432 7297 7460
rect 5960 7420 5966 7432
rect 7285 7429 7297 7432
rect 7331 7429 7343 7463
rect 8570 7460 8576 7472
rect 8531 7432 8576 7460
rect 7285 7423 7343 7429
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 12066 7460 12072 7472
rect 9798 7432 12072 7460
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 12618 7420 12624 7472
rect 12676 7420 12682 7472
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 13872 7432 14473 7460
rect 13872 7420 13878 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 15289 7463 15347 7469
rect 15289 7429 15301 7463
rect 15335 7460 15347 7463
rect 15378 7460 15384 7472
rect 15335 7432 15384 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 17405 7463 17463 7469
rect 17405 7429 17417 7463
rect 17451 7460 17463 7463
rect 18414 7460 18420 7472
rect 17451 7432 18420 7460
rect 17451 7429 17463 7432
rect 17405 7423 17463 7429
rect 18414 7420 18420 7432
rect 18472 7420 18478 7472
rect 19444 7469 19472 7500
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 22741 7531 22799 7537
rect 22741 7528 22753 7531
rect 21692 7500 22753 7528
rect 21692 7488 21698 7500
rect 22741 7497 22753 7500
rect 22787 7497 22799 7531
rect 22741 7491 22799 7497
rect 23014 7488 23020 7540
rect 23072 7528 23078 7540
rect 23385 7531 23443 7537
rect 23385 7528 23397 7531
rect 23072 7500 23397 7528
rect 23072 7488 23078 7500
rect 23385 7497 23397 7500
rect 23431 7497 23443 7531
rect 25222 7528 25228 7540
rect 25183 7500 25228 7528
rect 23385 7491 23443 7497
rect 25222 7488 25228 7500
rect 25280 7488 25286 7540
rect 19429 7463 19487 7469
rect 19429 7429 19441 7463
rect 19475 7429 19487 7463
rect 19429 7423 19487 7429
rect 19702 7420 19708 7472
rect 19760 7460 19766 7472
rect 20438 7460 20444 7472
rect 19760 7432 20444 7460
rect 19760 7420 19766 7432
rect 20438 7420 20444 7432
rect 20496 7420 20502 7472
rect 20622 7460 20628 7472
rect 20583 7432 20628 7460
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 20717 7463 20775 7469
rect 20717 7429 20729 7463
rect 20763 7460 20775 7463
rect 20990 7460 20996 7472
rect 20763 7432 20996 7460
rect 20763 7429 20775 7432
rect 20717 7423 20775 7429
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 21266 7420 21272 7472
rect 21324 7460 21330 7472
rect 22097 7463 22155 7469
rect 22097 7460 22109 7463
rect 21324 7432 22109 7460
rect 21324 7420 21330 7432
rect 22097 7429 22109 7432
rect 22143 7429 22155 7463
rect 22097 7423 22155 7429
rect 1394 7352 1400 7404
rect 1452 7392 1458 7404
rect 1765 7395 1823 7401
rect 1765 7392 1777 7395
rect 1452 7364 1777 7392
rect 1452 7352 1458 7364
rect 1765 7361 1777 7364
rect 1811 7361 1823 7395
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 1765 7355 1823 7361
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 4522 7392 4528 7404
rect 4483 7364 4528 7392
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5258 7392 5264 7404
rect 5215 7364 5264 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5810 7392 5816 7404
rect 5592 7364 5816 7392
rect 5592 7352 5598 7364
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 6546 7392 6552 7404
rect 6507 7364 6552 7392
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 8110 7392 8116 7404
rect 6696 7364 8116 7392
rect 6696 7352 6702 7364
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8297 7395 8355 7401
rect 8297 7392 8309 7395
rect 8220 7364 8309 7392
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4062 7324 4068 7336
rect 4019 7296 4068 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5132 7296 5917 7324
rect 5132 7284 5138 7296
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 8220 7324 8248 7364
rect 8297 7361 8309 7364
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10410 7392 10416 7404
rect 10100 7364 10416 7392
rect 10100 7352 10106 7364
rect 10410 7352 10416 7364
rect 10468 7392 10474 7404
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10468 7364 10609 7392
rect 10468 7352 10474 7364
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 10686 7352 10692 7404
rect 10744 7392 10750 7404
rect 14182 7392 14188 7404
rect 10744 7364 10789 7392
rect 14143 7364 14188 7392
rect 10744 7352 10750 7364
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 22002 7392 22008 7404
rect 21963 7364 22008 7392
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 23293 7395 23351 7401
rect 23293 7361 23305 7395
rect 23339 7392 23351 7395
rect 24210 7392 24216 7404
rect 23339 7364 24216 7392
rect 23339 7361 23351 7364
rect 23293 7355 23351 7361
rect 6972 7296 8248 7324
rect 6972 7284 6978 7296
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 11238 7324 11244 7336
rect 8628 7296 11244 7324
rect 8628 7284 8634 7296
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11664 7296 11897 7324
rect 11664 7284 11670 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 11885 7287 11943 7293
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7324 12219 7327
rect 14918 7324 14924 7336
rect 12207 7296 14924 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7324 15255 7327
rect 15286 7324 15292 7336
rect 15243 7296 15292 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 17310 7324 17316 7336
rect 17271 7296 17316 7324
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 17770 7324 17776 7336
rect 17731 7296 17776 7324
rect 17770 7284 17776 7296
rect 17828 7284 17834 7336
rect 18322 7284 18328 7336
rect 18380 7324 18386 7336
rect 19150 7324 19156 7336
rect 18380 7296 19156 7324
rect 18380 7284 18386 7296
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19337 7327 19395 7333
rect 19337 7293 19349 7327
rect 19383 7324 19395 7327
rect 19702 7324 19708 7336
rect 19383 7296 19708 7324
rect 19383 7293 19395 7296
rect 19337 7287 19395 7293
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 20254 7324 20260 7336
rect 19852 7296 20260 7324
rect 19852 7284 19858 7296
rect 20254 7284 20260 7296
rect 20312 7324 20318 7336
rect 20901 7327 20959 7333
rect 20901 7324 20913 7327
rect 20312 7296 20913 7324
rect 20312 7284 20318 7296
rect 20901 7293 20913 7296
rect 20947 7293 20959 7327
rect 20901 7287 20959 7293
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 22664 7324 22692 7355
rect 24210 7352 24216 7364
rect 24268 7352 24274 7404
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7392 24455 7395
rect 25038 7392 25044 7404
rect 24443 7364 25044 7392
rect 24443 7361 24455 7364
rect 24397 7355 24455 7361
rect 25038 7352 25044 7364
rect 25096 7352 25102 7404
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 21324 7296 22692 7324
rect 21324 7284 21330 7296
rect 23382 7284 23388 7336
rect 23440 7324 23446 7336
rect 23937 7327 23995 7333
rect 23937 7324 23949 7327
rect 23440 7296 23949 7324
rect 23440 7284 23446 7296
rect 23937 7293 23949 7296
rect 23983 7293 23995 7327
rect 24854 7324 24860 7336
rect 24815 7296 24860 7324
rect 23937 7287 23995 7293
rect 24854 7284 24860 7296
rect 24912 7324 24918 7336
rect 25424 7324 25452 7355
rect 24912 7296 25452 7324
rect 24912 7284 24918 7296
rect 4617 7259 4675 7265
rect 3804 7228 4108 7256
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 3804 7188 3832 7228
rect 1627 7160 3832 7188
rect 4080 7188 4108 7228
rect 4617 7225 4629 7259
rect 4663 7256 4675 7259
rect 15749 7259 15807 7265
rect 4663 7228 8432 7256
rect 4663 7225 4675 7228
rect 4617 7219 4675 7225
rect 4798 7188 4804 7200
rect 4080 7160 4804 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 8294 7188 8300 7200
rect 5040 7160 8300 7188
rect 5040 7148 5046 7160
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 8404 7188 8432 7228
rect 15749 7225 15761 7259
rect 15795 7256 15807 7259
rect 19058 7256 19064 7268
rect 15795 7228 19064 7256
rect 15795 7225 15807 7228
rect 15749 7219 15807 7225
rect 19058 7216 19064 7228
rect 19116 7216 19122 7268
rect 19889 7259 19947 7265
rect 19889 7256 19901 7259
rect 19306 7228 19901 7256
rect 9858 7188 9864 7200
rect 8404 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 12894 7188 12900 7200
rect 10091 7160 12900 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 16390 7188 16396 7200
rect 13679 7160 16396 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 18506 7188 18512 7200
rect 16540 7160 18512 7188
rect 16540 7148 16546 7160
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 18690 7148 18696 7200
rect 18748 7188 18754 7200
rect 19306 7188 19334 7228
rect 19889 7225 19901 7228
rect 19935 7256 19947 7259
rect 21818 7256 21824 7268
rect 19935 7228 21824 7256
rect 19935 7225 19947 7228
rect 19889 7219 19947 7225
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 18748 7160 19334 7188
rect 18748 7148 18754 7160
rect 23474 7148 23480 7200
rect 23532 7188 23538 7200
rect 24489 7191 24547 7197
rect 24489 7188 24501 7191
rect 23532 7160 24501 7188
rect 23532 7148 23538 7160
rect 24489 7157 24501 7160
rect 24535 7157 24547 7191
rect 24489 7151 24547 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1844 6987 1902 6993
rect 1844 6953 1856 6987
rect 1890 6984 1902 6987
rect 2038 6984 2044 6996
rect 1890 6956 2044 6984
rect 1890 6953 1902 6956
rect 1844 6947 1902 6953
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6162 6987 6220 6993
rect 6162 6984 6174 6987
rect 6052 6956 6174 6984
rect 6052 6944 6058 6956
rect 6162 6953 6174 6956
rect 6208 6953 6220 6987
rect 6162 6947 6220 6953
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7558 6984 7564 6996
rect 7248 6956 7564 6984
rect 7248 6944 7254 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 7708 6956 7753 6984
rect 7708 6944 7714 6956
rect 8202 6944 8208 6996
rect 8260 6984 8266 6996
rect 23198 6984 23204 6996
rect 8260 6956 23204 6984
rect 8260 6944 8266 6956
rect 23198 6944 23204 6956
rect 23256 6944 23262 6996
rect 8481 6919 8539 6925
rect 8481 6885 8493 6919
rect 8527 6916 8539 6919
rect 8527 6888 8616 6916
rect 8527 6885 8539 6888
rect 8481 6879 8539 6885
rect 3326 6848 3332 6860
rect 3239 6820 3332 6848
rect 3326 6808 3332 6820
rect 3384 6848 3390 6860
rect 3878 6848 3884 6860
rect 3384 6820 3884 6848
rect 3384 6808 3390 6820
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 4614 6848 4620 6860
rect 4264 6820 4620 6848
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 4264 6789 4292 6820
rect 4614 6808 4620 6820
rect 4672 6848 4678 6860
rect 6546 6848 6552 6860
rect 4672 6820 6552 6848
rect 4672 6808 4678 6820
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 5902 6780 5908 6792
rect 5863 6752 5908 6780
rect 4249 6743 4307 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 8202 6740 8208 6792
rect 8260 6782 8266 6792
rect 8381 6785 8439 6791
rect 8381 6782 8393 6785
rect 8260 6754 8393 6782
rect 8260 6740 8266 6754
rect 8381 6751 8393 6754
rect 8427 6751 8439 6785
rect 8588 6780 8616 6888
rect 8754 6876 8760 6928
rect 8812 6916 8818 6928
rect 9674 6916 9680 6928
rect 8812 6888 9680 6916
rect 8812 6876 8818 6888
rect 9674 6876 9680 6888
rect 9732 6876 9738 6928
rect 21634 6916 21640 6928
rect 12268 6888 21640 6916
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9766 6848 9772 6860
rect 8904 6820 9772 6848
rect 8904 6808 8910 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9030 6780 9036 6792
rect 8588 6752 9036 6780
rect 8381 6745 8439 6751
rect 9030 6740 9036 6752
rect 9088 6740 9094 6792
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9456 6752 9501 6780
rect 9456 6740 9462 6752
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9732 6752 10057 6780
rect 9732 6740 9738 6752
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 12268 6780 12296 6888
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 22112 6888 22508 6916
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 13998 6848 14004 6860
rect 13587 6820 14004 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14182 6848 14188 6860
rect 14108 6820 14188 6848
rect 11454 6752 12296 6780
rect 12345 6783 12403 6789
rect 10045 6743 10103 6749
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 12391 6752 13277 6780
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 13265 6749 13277 6752
rect 13311 6780 13323 6783
rect 14108 6780 14136 6820
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 14734 6848 14740 6860
rect 14415 6820 14740 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 15013 6851 15071 6857
rect 15013 6817 15025 6851
rect 15059 6848 15071 6851
rect 15286 6848 15292 6860
rect 15059 6820 15292 6848
rect 15059 6817 15071 6820
rect 15013 6811 15071 6817
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6848 15715 6851
rect 16482 6848 16488 6860
rect 15703 6820 16488 6848
rect 15703 6817 15715 6820
rect 15657 6811 15715 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16669 6851 16727 6857
rect 16669 6817 16681 6851
rect 16715 6848 16727 6851
rect 17126 6848 17132 6860
rect 16715 6820 17132 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 17310 6848 17316 6860
rect 17271 6820 17316 6848
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 19150 6848 19156 6860
rect 17696 6820 19156 6848
rect 14274 6780 14280 6792
rect 13311 6752 14136 6780
rect 14235 6752 14280 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 4614 6712 4620 6724
rect 3082 6684 4620 6712
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 4982 6712 4988 6724
rect 4943 6684 4988 6712
rect 4982 6672 4988 6684
rect 5040 6672 5046 6724
rect 8110 6712 8116 6724
rect 7406 6684 8116 6712
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 10318 6712 10324 6724
rect 10279 6684 10324 6712
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 12621 6715 12679 6721
rect 12621 6681 12633 6715
rect 12667 6712 12679 6715
rect 12710 6712 12716 6724
rect 12667 6684 12716 6712
rect 12667 6681 12679 6684
rect 12621 6675 12679 6681
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13814 6712 13820 6724
rect 12952 6684 13820 6712
rect 12952 6672 12958 6684
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 16761 6715 16819 6721
rect 15160 6684 15205 6712
rect 15160 6672 15166 6684
rect 16761 6681 16773 6715
rect 16807 6712 16819 6715
rect 17126 6712 17132 6724
rect 16807 6684 17132 6712
rect 16807 6681 16819 6684
rect 16761 6675 16819 6681
rect 17126 6672 17132 6684
rect 17184 6672 17190 6724
rect 17310 6672 17316 6724
rect 17368 6712 17374 6724
rect 17586 6712 17592 6724
rect 17368 6684 17592 6712
rect 17368 6672 17374 6684
rect 17586 6672 17592 6684
rect 17644 6672 17650 6724
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 9493 6647 9551 6653
rect 9493 6644 9505 6647
rect 7616 6616 9505 6644
rect 7616 6604 7622 6616
rect 9493 6613 9505 6616
rect 9539 6613 9551 6647
rect 9493 6607 9551 6613
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 11054 6644 11060 6656
rect 9640 6616 11060 6644
rect 9640 6604 9646 6616
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11330 6604 11336 6656
rect 11388 6644 11394 6656
rect 11793 6647 11851 6653
rect 11793 6644 11805 6647
rect 11388 6616 11805 6644
rect 11388 6604 11394 6616
rect 11793 6613 11805 6616
rect 11839 6613 11851 6647
rect 11793 6607 11851 6613
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 13354 6644 13360 6656
rect 11940 6616 13360 6644
rect 11940 6604 11946 6616
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 17696 6644 17724 6820
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 19521 6851 19579 6857
rect 19521 6848 19533 6851
rect 19352 6820 19533 6848
rect 19352 6792 19380 6820
rect 19521 6817 19533 6820
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 19886 6808 19892 6860
rect 19944 6848 19950 6860
rect 21361 6851 21419 6857
rect 19944 6820 21312 6848
rect 19944 6808 19950 6820
rect 19334 6740 19340 6792
rect 19392 6740 19398 6792
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6780 20223 6783
rect 20254 6780 20260 6792
rect 20211 6752 20260 6780
rect 20211 6749 20223 6752
rect 20165 6743 20223 6749
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21284 6780 21312 6820
rect 21361 6817 21373 6851
rect 21407 6848 21419 6851
rect 22112 6848 22140 6888
rect 22373 6851 22431 6857
rect 22373 6848 22385 6851
rect 21407 6820 22140 6848
rect 22204 6820 22385 6848
rect 21407 6817 21419 6820
rect 21361 6811 21419 6817
rect 22204 6780 22232 6820
rect 22373 6817 22385 6820
rect 22419 6817 22431 6851
rect 22480 6848 22508 6888
rect 23382 6848 23388 6860
rect 22480 6820 23244 6848
rect 23343 6820 23388 6848
rect 22373 6811 22431 6817
rect 21284 6752 22232 6780
rect 22281 6783 22339 6789
rect 21177 6743 21235 6749
rect 22281 6749 22293 6783
rect 22327 6780 22339 6783
rect 22646 6780 22652 6792
rect 22327 6752 22652 6780
rect 22327 6749 22339 6752
rect 22281 6743 22339 6749
rect 18141 6715 18199 6721
rect 18141 6681 18153 6715
rect 18187 6681 18199 6715
rect 18141 6675 18199 6681
rect 15252 6616 17724 6644
rect 18156 6644 18184 6675
rect 18230 6672 18236 6724
rect 18288 6712 18294 6724
rect 18288 6684 18333 6712
rect 18288 6672 18294 6684
rect 18506 6672 18512 6724
rect 18564 6712 18570 6724
rect 18785 6715 18843 6721
rect 18785 6712 18797 6715
rect 18564 6684 18797 6712
rect 18564 6672 18570 6684
rect 18785 6681 18797 6684
rect 18831 6681 18843 6715
rect 18785 6675 18843 6681
rect 18874 6672 18880 6724
rect 18932 6712 18938 6724
rect 19613 6715 19671 6721
rect 18932 6684 19564 6712
rect 18932 6672 18938 6684
rect 19334 6644 19340 6656
rect 18156 6616 19340 6644
rect 15252 6604 15258 6616
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19536 6644 19564 6684
rect 19613 6681 19625 6715
rect 19659 6712 19671 6715
rect 19702 6712 19708 6724
rect 19659 6684 19708 6712
rect 19659 6681 19671 6684
rect 19613 6675 19671 6681
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 21192 6712 21220 6743
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 23216 6780 23244 6820
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 23474 6780 23480 6792
rect 23216 6752 23480 6780
rect 23474 6740 23480 6752
rect 23532 6740 23538 6792
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 24581 6783 24639 6789
rect 23624 6752 23669 6780
rect 23624 6740 23630 6752
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24670 6780 24676 6792
rect 24627 6752 24676 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 21358 6712 21364 6724
rect 21192 6684 21364 6712
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 21174 6644 21180 6656
rect 19536 6616 21180 6644
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 21818 6644 21824 6656
rect 21731 6616 21824 6644
rect 21818 6604 21824 6616
rect 21876 6644 21882 6656
rect 22002 6644 22008 6656
rect 21876 6616 22008 6644
rect 21876 6604 21882 6616
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 24029 6647 24087 6653
rect 24029 6644 24041 6647
rect 22244 6616 24041 6644
rect 22244 6604 22250 6616
rect 24029 6613 24041 6616
rect 24075 6613 24087 6647
rect 24670 6644 24676 6656
rect 24631 6616 24676 6644
rect 24029 6607 24087 6613
rect 24670 6604 24676 6616
rect 24728 6604 24734 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 5902 6440 5908 6452
rect 4264 6412 5908 6440
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 4264 6313 4292 6412
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 11882 6440 11888 6452
rect 6748 6412 11888 6440
rect 6362 6372 6368 6384
rect 5750 6344 6368 6372
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3789 6307 3847 6313
rect 3789 6304 3801 6307
rect 3099 6276 3801 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3789 6273 3801 6276
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 2976 6236 3004 6267
rect 4525 6239 4583 6245
rect 2976 6208 4384 6236
rect 3605 6171 3663 6177
rect 3605 6168 3617 6171
rect 2746 6140 3617 6168
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 2314 6100 2320 6112
rect 1811 6072 2320 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2746 6100 2774 6140
rect 3605 6137 3617 6140
rect 3651 6137 3663 6171
rect 3605 6131 3663 6137
rect 2464 6072 2774 6100
rect 4356 6100 4384 6208
rect 4525 6205 4537 6239
rect 4571 6236 4583 6239
rect 6748 6236 6776 6412
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 17586 6440 17592 6452
rect 12360 6412 17592 6440
rect 7190 6372 7196 6384
rect 7151 6344 7196 6372
rect 7190 6332 7196 6344
rect 7248 6332 7254 6384
rect 9030 6372 9036 6384
rect 8418 6344 9036 6372
rect 9030 6332 9036 6344
rect 9088 6332 9094 6384
rect 9306 6372 9312 6384
rect 9140 6344 9312 6372
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 9140 6313 9168 6344
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9456 6344 9501 6372
rect 9456 6332 9462 6344
rect 9858 6332 9864 6384
rect 9916 6332 9922 6384
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 12360 6372 12388 6412
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 20622 6440 20628 6452
rect 17689 6412 20628 6440
rect 14185 6375 14243 6381
rect 14185 6372 14197 6375
rect 11480 6344 12388 6372
rect 13648 6344 14197 6372
rect 11480 6332 11486 6344
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 6880 6276 6929 6304
rect 6880 6264 6886 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 13078 6264 13084 6316
rect 13136 6264 13142 6316
rect 8202 6236 8208 6248
rect 4571 6208 6776 6236
rect 7024 6208 8208 6236
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 6546 6128 6552 6180
rect 6604 6168 6610 6180
rect 7024 6168 7052 6208
rect 8202 6196 8208 6208
rect 8260 6236 8266 6248
rect 9950 6236 9956 6248
rect 8260 6208 9956 6236
rect 8260 6196 8266 6208
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10870 6236 10876 6248
rect 10831 6208 10876 6236
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11238 6196 11244 6248
rect 11296 6236 11302 6248
rect 11606 6236 11612 6248
rect 11296 6208 11612 6236
rect 11296 6196 11302 6208
rect 11606 6196 11612 6208
rect 11664 6236 11670 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11664 6208 11713 6236
rect 11664 6196 11670 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6236 12035 6239
rect 12342 6236 12348 6248
rect 12023 6208 12348 6236
rect 12023 6205 12035 6208
rect 11977 6199 12035 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 13648 6168 13676 6344
rect 14185 6341 14197 6344
rect 14231 6341 14243 6375
rect 14185 6335 14243 6341
rect 14918 6332 14924 6384
rect 14976 6372 14982 6384
rect 15105 6375 15163 6381
rect 15105 6372 15117 6375
rect 14976 6344 15117 6372
rect 14976 6332 14982 6344
rect 15105 6341 15117 6344
rect 15151 6341 15163 6375
rect 15105 6335 15163 6341
rect 15749 6375 15807 6381
rect 15749 6341 15761 6375
rect 15795 6372 15807 6375
rect 17218 6372 17224 6384
rect 15795 6344 17224 6372
rect 15795 6341 15807 6344
rect 15749 6335 15807 6341
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 17689 6381 17717 6412
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20772 6412 21005 6440
rect 20772 6400 20778 6412
rect 20993 6409 21005 6412
rect 21039 6409 21051 6443
rect 20993 6403 21051 6409
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 22462 6440 22468 6452
rect 21232 6412 22468 6440
rect 21232 6400 21238 6412
rect 22462 6400 22468 6412
rect 22520 6400 22526 6452
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 22741 6443 22799 6449
rect 22741 6440 22753 6443
rect 22612 6412 22753 6440
rect 22612 6400 22618 6412
rect 22741 6409 22753 6412
rect 22787 6409 22799 6443
rect 22741 6403 22799 6409
rect 23566 6400 23572 6452
rect 23624 6440 23630 6452
rect 27157 6443 27215 6449
rect 27157 6440 27169 6443
rect 23624 6412 27169 6440
rect 23624 6400 23630 6412
rect 27157 6409 27169 6412
rect 27203 6409 27215 6443
rect 27157 6403 27215 6409
rect 30374 6400 30380 6452
rect 30432 6440 30438 6452
rect 32401 6443 32459 6449
rect 32401 6440 32413 6443
rect 30432 6412 32413 6440
rect 30432 6400 30438 6412
rect 32401 6409 32413 6412
rect 32447 6409 32459 6443
rect 38102 6440 38108 6452
rect 38063 6412 38108 6440
rect 32401 6403 32459 6409
rect 38102 6400 38108 6412
rect 38160 6400 38166 6452
rect 17681 6375 17739 6381
rect 17681 6341 17693 6375
rect 17727 6341 17739 6375
rect 18598 6372 18604 6384
rect 17681 6335 17739 6341
rect 18248 6344 18604 6372
rect 18248 6316 18276 6344
rect 18598 6332 18604 6344
rect 18656 6332 18662 6384
rect 18782 6372 18788 6384
rect 18743 6344 18788 6372
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 19794 6372 19800 6384
rect 19306 6344 19800 6372
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16853 6307 16911 6313
rect 16356 6276 16401 6304
rect 16356 6264 16362 6276
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 17310 6304 17316 6316
rect 16899 6276 17316 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18288 6276 18333 6304
rect 18288 6264 18294 6276
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18564 6276 18705 6304
rect 18564 6264 18570 6276
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 19306 6304 19334 6344
rect 19794 6332 19800 6344
rect 19852 6332 19858 6384
rect 19889 6375 19947 6381
rect 19889 6341 19901 6375
rect 19935 6372 19947 6375
rect 20530 6372 20536 6384
rect 19935 6344 20536 6372
rect 19935 6341 19947 6344
rect 19889 6335 19947 6341
rect 20530 6332 20536 6344
rect 20588 6332 20594 6384
rect 21450 6372 21456 6384
rect 20640 6344 21456 6372
rect 18739 6276 19334 6304
rect 20441 6307 20499 6313
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 20441 6273 20453 6307
rect 20487 6304 20499 6307
rect 20640 6304 20668 6344
rect 21450 6332 21456 6344
rect 21508 6332 21514 6384
rect 21910 6372 21916 6384
rect 21652 6344 21916 6372
rect 20487 6276 20668 6304
rect 20901 6307 20959 6313
rect 20487 6273 20499 6276
rect 20441 6267 20499 6273
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 21082 6304 21088 6316
rect 20947 6276 21088 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 21082 6264 21088 6276
rect 21140 6304 21146 6316
rect 21652 6304 21680 6344
rect 21910 6332 21916 6344
rect 21968 6332 21974 6384
rect 23385 6375 23443 6381
rect 23385 6372 23397 6375
rect 22572 6344 23397 6372
rect 21140 6276 21680 6304
rect 21140 6264 21146 6276
rect 21726 6264 21732 6316
rect 21784 6304 21790 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21784 6276 22017 6304
rect 21784 6264 21790 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22152 6276 22197 6304
rect 22152 6264 22158 6276
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 15194 6236 15200 6248
rect 14139 6208 15200 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 15657 6239 15715 6245
rect 15657 6205 15669 6239
rect 15703 6236 15715 6239
rect 16482 6236 16488 6248
rect 15703 6208 16488 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 16942 6236 16948 6248
rect 16903 6208 16948 6236
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6236 17647 6239
rect 18322 6236 18328 6248
rect 17635 6208 18328 6236
rect 17635 6205 17647 6208
rect 17589 6199 17647 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 18966 6196 18972 6248
rect 19024 6196 19030 6248
rect 19797 6239 19855 6245
rect 19797 6205 19809 6239
rect 19843 6236 19855 6239
rect 19843 6208 20576 6236
rect 19843 6205 19855 6208
rect 19797 6199 19855 6205
rect 6604 6140 7052 6168
rect 13280 6140 13676 6168
rect 18984 6168 19012 6196
rect 20548 6168 20576 6208
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 22572 6236 22600 6344
rect 23385 6341 23397 6344
rect 23431 6341 23443 6375
rect 23385 6335 23443 6341
rect 24394 6332 24400 6384
rect 24452 6372 24458 6384
rect 24673 6375 24731 6381
rect 24673 6372 24685 6375
rect 24452 6344 24685 6372
rect 24452 6332 24458 6344
rect 24673 6341 24685 6344
rect 24719 6341 24731 6375
rect 24673 6335 24731 6341
rect 22649 6307 22707 6313
rect 22649 6273 22661 6307
rect 22695 6304 22707 6307
rect 22922 6304 22928 6316
rect 22695 6276 22928 6304
rect 22695 6273 22707 6276
rect 22649 6267 22707 6273
rect 22922 6264 22928 6276
rect 22980 6264 22986 6316
rect 23290 6304 23296 6316
rect 23251 6276 23296 6304
rect 23290 6264 23296 6276
rect 23348 6264 23354 6316
rect 23934 6304 23940 6316
rect 23895 6276 23940 6304
rect 23934 6264 23940 6276
rect 23992 6264 23998 6316
rect 24581 6307 24639 6313
rect 24581 6273 24593 6307
rect 24627 6273 24639 6307
rect 24581 6267 24639 6273
rect 25317 6307 25375 6313
rect 25317 6273 25329 6307
rect 25363 6304 25375 6307
rect 26142 6304 26148 6316
rect 25363 6276 26004 6304
rect 26103 6276 26148 6304
rect 25363 6273 25375 6276
rect 25317 6267 25375 6273
rect 20680 6208 22600 6236
rect 20680 6196 20686 6208
rect 22830 6196 22836 6248
rect 22888 6236 22894 6248
rect 24596 6236 24624 6267
rect 22888 6208 24624 6236
rect 25976 6236 26004 6276
rect 26142 6264 26148 6276
rect 26200 6264 26206 6316
rect 26418 6264 26424 6316
rect 26476 6304 26482 6316
rect 27341 6307 27399 6313
rect 27341 6304 27353 6307
rect 26476 6276 27353 6304
rect 26476 6264 26482 6276
rect 27341 6273 27353 6276
rect 27387 6273 27399 6307
rect 27341 6267 27399 6273
rect 32309 6307 32367 6313
rect 32309 6273 32321 6307
rect 32355 6304 32367 6307
rect 34054 6304 34060 6316
rect 32355 6276 34060 6304
rect 32355 6273 32367 6276
rect 32309 6267 32367 6273
rect 34054 6264 34060 6276
rect 34112 6264 34118 6316
rect 38286 6304 38292 6316
rect 38247 6276 38292 6304
rect 38286 6264 38292 6276
rect 38344 6264 38350 6316
rect 28442 6236 28448 6248
rect 25976 6208 28448 6236
rect 22888 6196 22894 6208
rect 28442 6196 28448 6208
rect 28500 6196 28506 6248
rect 21818 6168 21824 6180
rect 18984 6140 20484 6168
rect 20548 6140 21824 6168
rect 6604 6128 6610 6140
rect 4890 6100 4896 6112
rect 4356 6072 4896 6100
rect 2464 6060 2470 6072
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 5994 6100 6000 6112
rect 5955 6072 6000 6100
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 10870 6100 10876 6112
rect 8711 6072 10876 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 13280 6100 13308 6140
rect 11112 6072 13308 6100
rect 11112 6060 11118 6072
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 13412 6072 13461 6100
rect 13412 6060 13418 6072
rect 13449 6069 13461 6072
rect 13495 6100 13507 6103
rect 16574 6100 16580 6112
rect 13495 6072 16580 6100
rect 13495 6069 13507 6072
rect 13449 6063 13507 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 18598 6100 18604 6112
rect 17276 6072 18604 6100
rect 17276 6060 17282 6072
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 19150 6060 19156 6112
rect 19208 6100 19214 6112
rect 20346 6100 20352 6112
rect 19208 6072 20352 6100
rect 19208 6060 19214 6072
rect 20346 6060 20352 6072
rect 20404 6060 20410 6112
rect 20456 6100 20484 6140
rect 21818 6128 21824 6140
rect 21876 6128 21882 6180
rect 24029 6171 24087 6177
rect 24029 6168 24041 6171
rect 21928 6140 24041 6168
rect 21928 6100 21956 6140
rect 24029 6137 24041 6140
rect 24075 6137 24087 6171
rect 24029 6131 24087 6137
rect 20456 6072 21956 6100
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 25409 6103 25467 6109
rect 25409 6100 25421 6103
rect 22060 6072 25421 6100
rect 22060 6060 22066 6072
rect 25409 6069 25421 6072
rect 25455 6069 25467 6103
rect 25409 6063 25467 6069
rect 25590 6060 25596 6112
rect 25648 6100 25654 6112
rect 25961 6103 26019 6109
rect 25961 6100 25973 6103
rect 25648 6072 25973 6100
rect 25648 6060 25654 6072
rect 25961 6069 25973 6072
rect 26007 6069 26019 6103
rect 25961 6063 26019 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 5905 5899 5963 5905
rect 3476 5868 5488 5896
rect 3476 5856 3482 5868
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1636 5732 1685 5760
rect 1636 5720 1642 5732
rect 1673 5729 1685 5732
rect 1719 5760 1731 5763
rect 2038 5760 2044 5772
rect 1719 5732 2044 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 2038 5720 2044 5732
rect 2096 5720 2102 5772
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5760 4215 5763
rect 4982 5760 4988 5772
rect 4203 5732 4988 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5460 5760 5488 5868
rect 5905 5865 5917 5899
rect 5951 5896 5963 5899
rect 6454 5896 6460 5908
rect 5951 5868 6460 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 8386 5896 8392 5908
rect 6564 5868 8392 5896
rect 5626 5788 5632 5840
rect 5684 5828 5690 5840
rect 6564 5828 6592 5868
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 11882 5896 11888 5908
rect 8619 5868 11888 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 20714 5896 20720 5908
rect 13136 5868 20720 5896
rect 13136 5856 13142 5868
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 21692 5868 23857 5896
rect 21692 5856 21698 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 24854 5896 24860 5908
rect 24815 5868 24860 5896
rect 23845 5859 23903 5865
rect 24854 5856 24860 5868
rect 24912 5856 24918 5908
rect 26418 5896 26424 5908
rect 26379 5868 26424 5896
rect 26418 5856 26424 5868
rect 26476 5856 26482 5908
rect 5684 5800 6592 5828
rect 5684 5788 5690 5800
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 10410 5828 10416 5840
rect 8168 5800 10416 5828
rect 8168 5788 8174 5800
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 10594 5828 10600 5840
rect 10555 5800 10600 5828
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 12989 5831 13047 5837
rect 10928 5800 11376 5828
rect 10928 5788 10934 5800
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 5460 5732 7113 5760
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 7101 5723 7159 5729
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 9861 5763 9919 5769
rect 9861 5760 9873 5763
rect 7248 5732 9873 5760
rect 7248 5720 7254 5732
rect 9861 5729 9873 5732
rect 9907 5729 9919 5763
rect 11238 5760 11244 5772
rect 11199 5732 11244 5760
rect 9861 5723 9919 5729
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 11348 5760 11376 5800
rect 12728 5800 12940 5828
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 11348 5732 11529 5760
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11606 5720 11612 5772
rect 11664 5760 11670 5772
rect 12728 5760 12756 5800
rect 11664 5732 12756 5760
rect 12912 5760 12940 5800
rect 12989 5797 13001 5831
rect 13035 5828 13047 5831
rect 13262 5828 13268 5840
rect 13035 5800 13268 5828
rect 13035 5797 13047 5800
rect 12989 5791 13047 5797
rect 13262 5788 13268 5800
rect 13320 5788 13326 5840
rect 17126 5788 17132 5840
rect 17184 5828 17190 5840
rect 18598 5828 18604 5840
rect 17184 5800 18604 5828
rect 17184 5788 17190 5800
rect 18598 5788 18604 5800
rect 18656 5788 18662 5840
rect 19426 5788 19432 5840
rect 19484 5828 19490 5840
rect 19797 5831 19855 5837
rect 19797 5828 19809 5831
rect 19484 5800 19809 5828
rect 19484 5788 19490 5800
rect 19797 5797 19809 5800
rect 19843 5797 19855 5831
rect 19797 5791 19855 5797
rect 20254 5788 20260 5840
rect 20312 5828 20318 5840
rect 21913 5831 21971 5837
rect 21913 5828 21925 5831
rect 20312 5800 21925 5828
rect 20312 5788 20318 5800
rect 21913 5797 21925 5800
rect 21959 5797 21971 5831
rect 23201 5831 23259 5837
rect 23201 5828 23213 5831
rect 21913 5791 21971 5797
rect 22066 5800 23213 5828
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 12912 5732 14289 5760
rect 11664 5720 11670 5732
rect 14277 5729 14289 5732
rect 14323 5760 14335 5763
rect 14642 5760 14648 5772
rect 14323 5732 14648 5760
rect 14323 5729 14335 5732
rect 14277 5723 14335 5729
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 18012 5732 18245 5760
rect 18012 5720 18018 5732
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 6822 5692 6828 5704
rect 6783 5664 6828 5692
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 10134 5692 10140 5704
rect 8628 5664 10140 5692
rect 8628 5652 8634 5664
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5692 10563 5695
rect 10594 5692 10600 5704
rect 10551 5664 10600 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 16669 5695 16727 5701
rect 13596 5664 13641 5692
rect 13596 5652 13602 5664
rect 16669 5661 16681 5695
rect 16715 5692 16727 5695
rect 16758 5692 16764 5704
rect 16715 5664 16764 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 18248 5692 18276 5723
rect 18506 5720 18512 5772
rect 18564 5760 18570 5772
rect 20456 5769 20668 5772
rect 20456 5763 20683 5769
rect 20456 5760 20637 5763
rect 18564 5744 20637 5760
rect 18564 5732 20484 5744
rect 18564 5720 18570 5732
rect 20625 5729 20637 5744
rect 20671 5729 20683 5763
rect 20625 5723 20683 5729
rect 20898 5720 20904 5772
rect 20956 5760 20962 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20956 5732 21281 5760
rect 20956 5720 20962 5732
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 18322 5692 18328 5704
rect 18248 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 18748 5664 19441 5692
rect 18748 5652 18754 5664
rect 19429 5661 19441 5664
rect 19475 5692 19487 5695
rect 19518 5692 19524 5704
rect 19475 5664 19524 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 1949 5627 2007 5633
rect 1949 5593 1961 5627
rect 1995 5593 2007 5627
rect 4433 5627 4491 5633
rect 3174 5596 4384 5624
rect 1949 5587 2007 5593
rect 1964 5556 1992 5587
rect 3326 5556 3332 5568
rect 1964 5528 3332 5556
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 4356 5556 4384 5596
rect 4433 5593 4445 5627
rect 4479 5624 4491 5627
rect 4522 5624 4528 5636
rect 4479 5596 4528 5624
rect 4479 5593 4491 5596
rect 4433 5587 4491 5593
rect 4522 5584 4528 5596
rect 4580 5584 4586 5636
rect 6840 5624 6868 5652
rect 7190 5624 7196 5636
rect 6840 5596 7196 5624
rect 7190 5584 7196 5596
rect 7248 5584 7254 5636
rect 7558 5584 7564 5636
rect 7616 5584 7622 5636
rect 9125 5627 9183 5633
rect 9125 5593 9137 5627
rect 9171 5624 9183 5627
rect 9766 5624 9772 5636
rect 9171 5596 9772 5624
rect 9171 5593 9183 5596
rect 9125 5587 9183 5593
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 14458 5624 14464 5636
rect 11624 5596 12006 5624
rect 12820 5596 14464 5624
rect 8110 5556 8116 5568
rect 3476 5528 3521 5556
rect 4356 5528 8116 5556
rect 3476 5516 3482 5528
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8386 5516 8392 5568
rect 8444 5556 8450 5568
rect 11624 5556 11652 5596
rect 8444 5528 11652 5556
rect 8444 5516 8450 5528
rect 11882 5516 11888 5568
rect 11940 5556 11946 5568
rect 12820 5556 12848 5596
rect 14458 5584 14464 5596
rect 14516 5624 14522 5636
rect 14553 5627 14611 5633
rect 14553 5624 14565 5627
rect 14516 5596 14565 5624
rect 14516 5584 14522 5596
rect 14553 5593 14565 5596
rect 14599 5593 14611 5627
rect 14553 5587 14611 5593
rect 15010 5584 15016 5636
rect 15068 5584 15074 5636
rect 15930 5624 15936 5636
rect 15856 5596 15936 5624
rect 11940 5528 12848 5556
rect 13633 5559 13691 5565
rect 11940 5516 11946 5528
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 15856 5556 15884 5596
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 17402 5624 17408 5636
rect 17363 5596 17408 5624
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 17497 5627 17555 5633
rect 17497 5593 17509 5627
rect 17543 5624 17555 5627
rect 18506 5624 18512 5636
rect 17543 5596 18512 5624
rect 17543 5593 17555 5596
rect 17497 5587 17555 5593
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 19628 5624 19656 5655
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20533 5695 20591 5701
rect 20533 5692 20545 5695
rect 20404 5664 20545 5692
rect 20404 5652 20410 5664
rect 20533 5661 20545 5664
rect 20579 5692 20591 5695
rect 21082 5692 21088 5704
rect 20579 5664 21088 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 21082 5652 21088 5664
rect 21140 5652 21146 5704
rect 21177 5695 21235 5701
rect 21177 5661 21189 5695
rect 21223 5692 21235 5695
rect 21542 5692 21548 5704
rect 21223 5664 21548 5692
rect 21223 5661 21235 5664
rect 21177 5655 21235 5661
rect 21542 5652 21548 5664
rect 21600 5652 21606 5704
rect 21726 5652 21732 5704
rect 21784 5692 21790 5704
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 21784 5664 21833 5692
rect 21784 5652 21790 5664
rect 21821 5661 21833 5664
rect 21867 5661 21879 5695
rect 21821 5655 21879 5661
rect 22066 5624 22094 5800
rect 23201 5797 23213 5800
rect 23247 5797 23259 5831
rect 23201 5791 23259 5797
rect 23658 5788 23664 5840
rect 23716 5828 23722 5840
rect 24489 5831 24547 5837
rect 24489 5828 24501 5831
rect 23716 5800 24501 5828
rect 23716 5788 23722 5800
rect 24489 5797 24501 5800
rect 24535 5797 24547 5831
rect 24489 5791 24547 5797
rect 24872 5760 24900 5856
rect 25038 5788 25044 5840
rect 25096 5828 25102 5840
rect 25096 5800 25544 5828
rect 25096 5788 25102 5800
rect 24872 5732 25452 5760
rect 22462 5692 22468 5704
rect 22423 5664 22468 5692
rect 22462 5652 22468 5664
rect 22520 5652 22526 5704
rect 23106 5692 23112 5704
rect 23067 5664 23112 5692
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 25424 5701 25452 5732
rect 23753 5695 23811 5701
rect 23753 5661 23765 5695
rect 23799 5661 23811 5695
rect 23753 5655 23811 5661
rect 24397 5695 24455 5701
rect 24397 5661 24409 5695
rect 24443 5692 24455 5695
rect 25409 5695 25467 5701
rect 24443 5664 25268 5692
rect 24443 5661 24455 5664
rect 24397 5655 24455 5661
rect 23768 5624 23796 5655
rect 19628 5596 22094 5624
rect 22296 5596 23796 5624
rect 16022 5556 16028 5568
rect 13679 5528 15884 5556
rect 15983 5528 16028 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 16114 5516 16120 5568
rect 16172 5556 16178 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 16172 5528 16681 5556
rect 16172 5516 16178 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 16669 5519 16727 5525
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 21450 5556 21456 5568
rect 16816 5528 21456 5556
rect 16816 5516 16822 5528
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 21818 5516 21824 5568
rect 21876 5556 21882 5568
rect 22296 5556 22324 5596
rect 21876 5528 22324 5556
rect 21876 5516 21882 5528
rect 22370 5516 22376 5568
rect 22428 5556 22434 5568
rect 25240 5565 25268 5664
rect 25409 5661 25421 5695
rect 25455 5661 25467 5695
rect 25516 5692 25544 5800
rect 26605 5695 26663 5701
rect 26605 5692 26617 5695
rect 25516 5664 26617 5692
rect 25409 5655 25467 5661
rect 26605 5661 26617 5664
rect 26651 5661 26663 5695
rect 26605 5655 26663 5661
rect 22557 5559 22615 5565
rect 22557 5556 22569 5559
rect 22428 5528 22569 5556
rect 22428 5516 22434 5528
rect 22557 5525 22569 5528
rect 22603 5525 22615 5559
rect 22557 5519 22615 5525
rect 25225 5559 25283 5565
rect 25225 5525 25237 5559
rect 25271 5525 25283 5559
rect 25225 5519 25283 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 6822 5352 6828 5364
rect 4264 5324 6828 5352
rect 3878 5284 3884 5296
rect 3542 5256 3884 5284
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 4264 5225 4292 5324
rect 6822 5312 6828 5324
rect 6880 5352 6886 5364
rect 6880 5324 7144 5352
rect 6880 5312 6886 5324
rect 4430 5244 4436 5296
rect 4488 5284 4494 5296
rect 4525 5287 4583 5293
rect 4525 5284 4537 5287
rect 4488 5256 4537 5284
rect 4488 5244 4494 5256
rect 4525 5253 4537 5256
rect 4571 5253 4583 5287
rect 4525 5247 4583 5253
rect 4614 5244 4620 5296
rect 4672 5284 4678 5296
rect 4672 5256 5014 5284
rect 4672 5244 4678 5256
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 6546 5216 6552 5228
rect 6507 5188 6552 5216
rect 4249 5179 4307 5185
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 7116 5216 7144 5324
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 17586 5352 17592 5364
rect 9824 5324 13952 5352
rect 9824 5312 9830 5324
rect 9950 5284 9956 5296
rect 9416 5256 9956 5284
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 7116 5188 7205 5216
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 9416 5216 9444 5256
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 13924 5293 13952 5324
rect 15488 5324 17592 5352
rect 13909 5287 13967 5293
rect 13909 5253 13921 5287
rect 13955 5253 13967 5287
rect 14642 5284 14648 5296
rect 14603 5256 14648 5284
rect 13909 5247 13967 5253
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 9324 5188 9444 5216
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2682 5148 2688 5160
rect 2363 5120 2688 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3789 5151 3847 5157
rect 3789 5117 3801 5151
rect 3835 5148 3847 5151
rect 5166 5148 5172 5160
rect 3835 5120 5172 5148
rect 3835 5117 3847 5120
rect 3789 5111 3847 5117
rect 5166 5108 5172 5120
rect 5224 5148 5230 5160
rect 6270 5148 6276 5160
rect 5224 5120 6276 5148
rect 5224 5108 5230 5120
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6638 5108 6644 5160
rect 6696 5108 6702 5160
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 7834 5148 7840 5160
rect 7515 5120 7840 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 5718 5040 5724 5092
rect 5776 5080 5782 5092
rect 5997 5083 6055 5089
rect 5997 5080 6009 5083
rect 5776 5052 6009 5080
rect 5776 5040 5782 5052
rect 5997 5049 6009 5052
rect 6043 5080 6055 5083
rect 6656 5080 6684 5108
rect 9324 5080 9352 5188
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 15488 5216 15516 5324
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 20622 5352 20628 5364
rect 18340 5324 20628 5352
rect 15749 5287 15807 5293
rect 15749 5253 15761 5287
rect 15795 5284 15807 5287
rect 17313 5287 17371 5293
rect 15795 5256 17080 5284
rect 15795 5253 15807 5256
rect 15749 5247 15807 5253
rect 11296 5188 11744 5216
rect 13110 5188 15516 5216
rect 16301 5219 16359 5225
rect 11296 5176 11302 5188
rect 11716 5160 11744 5188
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16758 5216 16764 5228
rect 16347 5188 16764 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5148 9735 5151
rect 11698 5148 11704 5160
rect 9723 5120 11560 5148
rect 11659 5120 11704 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 6043 5052 6684 5080
rect 8864 5052 9352 5080
rect 6043 5049 6055 5052
rect 5997 5043 6055 5049
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 5258 5012 5264 5024
rect 4580 4984 5264 5012
rect 4580 4972 4586 4984
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 8864 5012 8892 5052
rect 6687 4984 8892 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 9416 5012 9444 5111
rect 11146 5080 11152 5092
rect 11107 5052 11152 5080
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 9674 5012 9680 5024
rect 8996 4984 9041 5012
rect 9416 4984 9680 5012
rect 8996 4972 9002 4984
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 11532 5012 11560 5120
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 15657 5151 15715 5157
rect 12023 5120 15608 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 15580 5080 15608 5120
rect 15657 5117 15669 5151
rect 15703 5148 15715 5151
rect 15838 5148 15844 5160
rect 15703 5120 15844 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 15930 5080 15936 5092
rect 15580 5052 15936 5080
rect 15930 5040 15936 5052
rect 15988 5040 15994 5092
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 17052 5080 17080 5256
rect 17313 5253 17325 5287
rect 17359 5284 17371 5287
rect 18340 5284 18368 5324
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 20916 5324 24685 5352
rect 18506 5284 18512 5296
rect 17359 5256 18368 5284
rect 18467 5256 18512 5284
rect 17359 5253 17371 5256
rect 17313 5247 17371 5253
rect 18506 5244 18512 5256
rect 18564 5244 18570 5296
rect 18690 5244 18696 5296
rect 18748 5284 18754 5296
rect 19058 5284 19064 5296
rect 18748 5256 19064 5284
rect 18748 5244 18754 5256
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 19150 5244 19156 5296
rect 19208 5284 19214 5296
rect 19702 5284 19708 5296
rect 19208 5256 19708 5284
rect 19208 5244 19214 5256
rect 19702 5244 19708 5256
rect 19760 5244 19766 5296
rect 19797 5287 19855 5293
rect 19797 5253 19809 5287
rect 19843 5284 19855 5287
rect 20806 5284 20812 5296
rect 19843 5256 20392 5284
rect 19843 5253 19855 5256
rect 19797 5247 19855 5253
rect 20364 5216 20392 5256
rect 20548 5256 20812 5284
rect 20438 5216 20444 5228
rect 20364 5188 20444 5216
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 17218 5148 17224 5160
rect 17179 5120 17224 5148
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 18417 5151 18475 5157
rect 17696 5120 18368 5148
rect 17696 5080 17724 5120
rect 16632 5052 16988 5080
rect 17052 5052 17724 5080
rect 16632 5040 16638 5052
rect 12158 5012 12164 5024
rect 11532 4984 12164 5012
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 13449 5015 13507 5021
rect 13449 5012 13461 5015
rect 13412 4984 13461 5012
rect 13412 4972 13418 4984
rect 13449 4981 13461 4984
rect 13495 4981 13507 5015
rect 13449 4975 13507 4981
rect 15286 4972 15292 5024
rect 15344 5012 15350 5024
rect 16850 5012 16856 5024
rect 15344 4984 16856 5012
rect 15344 4972 15350 4984
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 16960 5012 16988 5052
rect 17770 5040 17776 5092
rect 17828 5080 17834 5092
rect 18340 5080 18368 5120
rect 18417 5117 18429 5151
rect 18463 5148 18475 5151
rect 19426 5148 19432 5160
rect 18463 5120 19432 5148
rect 18463 5117 18475 5120
rect 18417 5111 18475 5117
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5148 19763 5151
rect 19886 5148 19892 5160
rect 19751 5120 19892 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 20349 5151 20407 5157
rect 20349 5148 20361 5151
rect 20036 5120 20361 5148
rect 20036 5108 20042 5120
rect 20349 5117 20361 5120
rect 20395 5148 20407 5151
rect 20548 5148 20576 5256
rect 20806 5244 20812 5256
rect 20864 5244 20870 5296
rect 20714 5176 20720 5228
rect 20772 5216 20778 5228
rect 20916 5216 20944 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 24673 5315 24731 5321
rect 21082 5244 21088 5296
rect 21140 5284 21146 5296
rect 21140 5256 21220 5284
rect 21140 5244 21146 5256
rect 20772 5188 20944 5216
rect 21077 5209 21135 5215
rect 20772 5176 20778 5188
rect 21077 5175 21089 5209
rect 21123 5200 21135 5209
rect 21192 5200 21220 5256
rect 22278 5244 22284 5296
rect 22336 5284 22342 5296
rect 22336 5256 23336 5284
rect 22336 5244 22342 5256
rect 21123 5175 21220 5200
rect 21266 5176 21272 5228
rect 21324 5216 21330 5228
rect 22462 5216 22468 5228
rect 21324 5188 22468 5216
rect 21324 5176 21330 5188
rect 22462 5176 22468 5188
rect 22520 5176 22526 5228
rect 22646 5216 22652 5228
rect 22607 5188 22652 5216
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 23308 5225 23336 5256
rect 23293 5219 23351 5225
rect 23293 5185 23305 5219
rect 23339 5185 23351 5219
rect 23293 5179 23351 5185
rect 23382 5176 23388 5228
rect 23440 5216 23446 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23440 5188 23949 5216
rect 23440 5176 23446 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24026 5176 24032 5228
rect 24084 5216 24090 5228
rect 24581 5219 24639 5225
rect 24581 5216 24593 5219
rect 24084 5188 24593 5216
rect 24084 5176 24090 5188
rect 24581 5185 24593 5188
rect 24627 5185 24639 5219
rect 24581 5179 24639 5185
rect 21077 5172 21220 5175
rect 21077 5169 21135 5172
rect 20395 5120 20576 5148
rect 20395 5117 20407 5120
rect 20349 5111 20407 5117
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 22005 5151 22063 5157
rect 22005 5148 22017 5151
rect 20864 5136 21036 5148
rect 21284 5136 22017 5148
rect 20864 5120 22017 5136
rect 20864 5108 20870 5120
rect 21008 5108 21312 5120
rect 22005 5117 22017 5120
rect 22051 5117 22063 5151
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 22005 5111 22063 5117
rect 22112 5120 22753 5148
rect 18874 5080 18880 5092
rect 17828 5052 17873 5080
rect 18340 5052 18880 5080
rect 17828 5040 17834 5052
rect 18874 5040 18880 5052
rect 18932 5040 18938 5092
rect 22112 5080 22140 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 24596 5148 24624 5179
rect 24946 5176 24952 5228
rect 25004 5216 25010 5228
rect 25409 5219 25467 5225
rect 25409 5216 25421 5219
rect 25004 5188 25421 5216
rect 25004 5176 25010 5188
rect 25409 5185 25421 5188
rect 25455 5185 25467 5219
rect 38010 5216 38016 5228
rect 37971 5188 38016 5216
rect 25409 5179 25467 5185
rect 38010 5176 38016 5188
rect 38068 5176 38074 5228
rect 24596 5120 25452 5148
rect 22741 5111 22799 5117
rect 25424 5092 25452 5120
rect 23385 5083 23443 5089
rect 23385 5080 23397 5083
rect 19812 5052 22140 5080
rect 22664 5052 23397 5080
rect 19812 5012 19840 5052
rect 16960 4984 19840 5012
rect 19886 4972 19892 5024
rect 19944 5012 19950 5024
rect 20622 5012 20628 5024
rect 19944 4984 20628 5012
rect 19944 4972 19950 4984
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 21174 5012 21180 5024
rect 21135 4984 21180 5012
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 21266 4972 21272 5024
rect 21324 5012 21330 5024
rect 22664 5012 22692 5052
rect 23385 5049 23397 5052
rect 23431 5049 23443 5083
rect 23385 5043 23443 5049
rect 23474 5040 23480 5092
rect 23532 5080 23538 5092
rect 23532 5052 24164 5080
rect 23532 5040 23538 5052
rect 21324 4984 22692 5012
rect 21324 4972 21330 4984
rect 22830 4972 22836 5024
rect 22888 5012 22894 5024
rect 24029 5015 24087 5021
rect 24029 5012 24041 5015
rect 22888 4984 24041 5012
rect 22888 4972 22894 4984
rect 24029 4981 24041 4984
rect 24075 4981 24087 5015
rect 24136 5012 24164 5052
rect 25406 5040 25412 5092
rect 25464 5040 25470 5092
rect 25225 5015 25283 5021
rect 25225 5012 25237 5015
rect 24136 4984 25237 5012
rect 24029 4975 24087 4981
rect 25225 4981 25237 4984
rect 25271 4981 25283 5015
rect 38194 5012 38200 5024
rect 38155 4984 38200 5012
rect 25225 4975 25283 4981
rect 38194 4972 38200 4984
rect 38252 4972 38258 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1844 4811 1902 4817
rect 1844 4777 1856 4811
rect 1890 4808 1902 4811
rect 3418 4808 3424 4820
rect 1890 4780 3424 4808
rect 1890 4777 1902 4780
rect 1844 4771 1902 4777
rect 3418 4768 3424 4780
rect 3476 4808 3482 4820
rect 4522 4808 4528 4820
rect 3476 4780 4528 4808
rect 3476 4768 3482 4780
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 5408 4780 7849 4808
rect 5408 4768 5414 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 10042 4808 10048 4820
rect 8444 4780 10048 4808
rect 8444 4768 8450 4780
rect 10042 4768 10048 4780
rect 10100 4808 10106 4820
rect 10686 4808 10692 4820
rect 10100 4780 10692 4808
rect 10100 4768 10106 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11320 4811 11378 4817
rect 11320 4777 11332 4811
rect 11366 4808 11378 4811
rect 12526 4808 12532 4820
rect 11366 4780 12532 4808
rect 11366 4777 11378 4780
rect 11320 4771 11378 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12805 4811 12863 4817
rect 12805 4777 12817 4811
rect 12851 4808 12863 4811
rect 12894 4808 12900 4820
rect 12851 4780 12900 4808
rect 12851 4777 12863 4780
rect 12805 4771 12863 4777
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 3602 4740 3608 4752
rect 3375 4712 3608 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 3602 4700 3608 4712
rect 3660 4700 3666 4752
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 6641 4743 6699 4749
rect 4764 4712 5028 4740
rect 4764 4700 4770 4712
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4672 1639 4675
rect 1946 4672 1952 4684
rect 1627 4644 1952 4672
rect 1627 4641 1639 4644
rect 1581 4635 1639 4641
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 3418 4632 3424 4684
rect 3476 4672 3482 4684
rect 3694 4672 3700 4684
rect 3476 4644 3700 4672
rect 3476 4632 3482 4644
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5000 4672 5028 4712
rect 6641 4709 6653 4743
rect 6687 4740 6699 4743
rect 6687 4712 8892 4740
rect 6687 4709 6699 4712
rect 6641 4703 6699 4709
rect 8481 4675 8539 4681
rect 8481 4672 8493 4675
rect 5000 4644 8493 4672
rect 8481 4641 8493 4644
rect 8527 4641 8539 4675
rect 8481 4635 8539 4641
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4706 4604 4712 4616
rect 4479 4576 4712 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7742 4604 7748 4616
rect 7064 4576 7748 4604
rect 7064 4564 7070 4576
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 8386 4604 8392 4616
rect 7892 4576 8392 4604
rect 7892 4564 7898 4576
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8864 4604 8892 4712
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 12820 4740 12848 4771
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13504 4780 13645 4808
rect 13504 4768 13510 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 14918 4768 14924 4820
rect 14976 4808 14982 4820
rect 17678 4808 17684 4820
rect 14976 4780 17684 4808
rect 14976 4768 14982 4780
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18138 4768 18144 4820
rect 18196 4808 18202 4820
rect 18509 4811 18567 4817
rect 18509 4808 18521 4811
rect 18196 4780 18521 4808
rect 18196 4768 18202 4780
rect 18509 4777 18521 4780
rect 18555 4777 18567 4811
rect 18509 4771 18567 4777
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 18932 4780 19472 4808
rect 18932 4768 18938 4780
rect 19334 4740 19340 4752
rect 12492 4712 12848 4740
rect 15764 4712 19340 4740
rect 12492 4700 12498 4712
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 10318 4672 10324 4684
rect 8996 4644 10324 4672
rect 8996 4632 9002 4644
rect 10318 4632 10324 4644
rect 10376 4672 10382 4684
rect 11974 4672 11980 4684
rect 10376 4644 11980 4672
rect 10376 4632 10382 4644
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 14240 4644 14289 4672
rect 14240 4632 14246 4644
rect 14277 4641 14289 4644
rect 14323 4672 14335 4675
rect 14642 4672 14648 4684
rect 14323 4644 14648 4672
rect 14323 4641 14335 4644
rect 14277 4635 14335 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 9677 4607 9735 4613
rect 8864 4576 9628 4604
rect 3694 4536 3700 4548
rect 3082 4508 3700 4536
rect 3694 4496 3700 4508
rect 3752 4496 3758 4548
rect 5166 4496 5172 4548
rect 5224 4536 5230 4548
rect 5224 4508 5269 4536
rect 5224 4496 5230 4508
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 9600 4536 9628 4576
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 9766 4604 9772 4616
rect 9723 4576 9772 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 10962 4604 10968 4616
rect 10551 4576 10968 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 10962 4564 10968 4576
rect 11020 4604 11026 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 11020 4576 11069 4604
rect 11020 4564 11026 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 14090 4604 14096 4616
rect 13587 4576 14096 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 15764 4604 15792 4712
rect 19334 4700 19340 4712
rect 19392 4700 19398 4752
rect 19444 4740 19472 4780
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19576 4780 19809 4808
rect 19576 4768 19582 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 19886 4768 19892 4820
rect 19944 4808 19950 4820
rect 20346 4808 20352 4820
rect 19944 4780 20352 4808
rect 19944 4768 19950 4780
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 20530 4808 20536 4820
rect 20491 4780 20536 4808
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 21269 4811 21327 4817
rect 21269 4808 21281 4811
rect 20640 4780 21281 4808
rect 20640 4740 20668 4780
rect 21269 4777 21281 4780
rect 21315 4777 21327 4811
rect 21269 4771 21327 4777
rect 21358 4768 21364 4820
rect 21416 4808 21422 4820
rect 23106 4808 23112 4820
rect 21416 4780 23112 4808
rect 21416 4768 21422 4780
rect 23106 4768 23112 4780
rect 23164 4768 23170 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 24486 4808 24492 4820
rect 23256 4780 23301 4808
rect 23400 4780 24492 4808
rect 23256 4768 23262 4780
rect 19444 4712 20668 4740
rect 22002 4700 22008 4752
rect 22060 4740 22066 4752
rect 23400 4740 23428 4780
rect 24486 4768 24492 4780
rect 24544 4768 24550 4820
rect 28166 4808 28172 4820
rect 24596 4780 26096 4808
rect 28127 4780 28172 4808
rect 22060 4712 23428 4740
rect 22060 4700 22066 4712
rect 16942 4672 16948 4684
rect 16903 4644 16948 4672
rect 16942 4632 16948 4644
rect 17000 4632 17006 4684
rect 17402 4632 17408 4684
rect 17460 4672 17466 4684
rect 17954 4672 17960 4684
rect 17460 4644 17816 4672
rect 17915 4644 17960 4672
rect 17460 4632 17466 4644
rect 15686 4576 15792 4604
rect 16574 4564 16580 4616
rect 16632 4564 16638 4616
rect 17788 4604 17816 4644
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 19426 4672 19432 4684
rect 18104 4644 18460 4672
rect 19387 4644 19432 4672
rect 18104 4632 18110 4644
rect 18432 4613 18460 4644
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 20162 4672 20168 4684
rect 19659 4644 20168 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 21266 4672 21272 4684
rect 20272 4644 21272 4672
rect 18417 4607 18475 4613
rect 17788 4576 18184 4604
rect 11422 4536 11428 4548
rect 5500 4508 5658 4536
rect 6472 4508 8064 4536
rect 9600 4508 11428 4536
rect 5500 4496 5506 4508
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 4982 4468 4988 4480
rect 4295 4440 4988 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 6472 4468 6500 4508
rect 5316 4440 6500 4468
rect 5316 4428 5322 4440
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 7926 4468 7932 4480
rect 6972 4440 7932 4468
rect 6972 4428 6978 4440
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8036 4468 8064 4508
rect 11422 4496 11428 4508
rect 11480 4496 11486 4548
rect 14274 4536 14280 4548
rect 12558 4508 14280 4536
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 14550 4536 14556 4548
rect 14511 4508 14556 4536
rect 14550 4496 14556 4508
rect 14608 4496 14614 4548
rect 16592 4536 16620 4564
rect 17030 4539 17088 4545
rect 17030 4536 17042 4539
rect 16592 4508 17042 4536
rect 17030 4505 17042 4508
rect 17076 4505 17088 4539
rect 18156 4536 18184 4576
rect 18417 4573 18429 4607
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 20272 4604 20300 4644
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 23382 4672 23388 4684
rect 22066 4644 23388 4672
rect 18656 4576 20300 4604
rect 18656 4564 18662 4576
rect 20346 4564 20352 4616
rect 20404 4604 20410 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20404 4576 20729 4604
rect 20404 4564 20410 4576
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 21177 4607 21235 4613
rect 21177 4604 21189 4607
rect 20717 4567 20775 4573
rect 20824 4576 21189 4604
rect 20530 4536 20536 4548
rect 18156 4508 20536 4536
rect 17030 4499 17088 4505
rect 20530 4496 20536 4508
rect 20588 4536 20594 4548
rect 20824 4536 20852 4576
rect 21177 4573 21189 4576
rect 21223 4573 21235 4607
rect 21177 4567 21235 4573
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4604 21879 4607
rect 22066 4604 22094 4644
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 24596 4672 24624 4780
rect 24854 4700 24860 4752
rect 24912 4740 24918 4752
rect 25869 4743 25927 4749
rect 25869 4740 25881 4743
rect 24912 4712 25881 4740
rect 24912 4700 24918 4712
rect 25869 4709 25881 4712
rect 25915 4709 25927 4743
rect 25869 4703 25927 4709
rect 23492 4644 24624 4672
rect 22462 4604 22468 4616
rect 21867 4576 22094 4604
rect 22423 4576 22468 4604
rect 21867 4573 21879 4576
rect 21821 4567 21879 4573
rect 22462 4564 22468 4576
rect 22520 4564 22526 4616
rect 23106 4604 23112 4616
rect 23067 4576 23112 4604
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 23290 4564 23296 4616
rect 23348 4604 23354 4616
rect 23492 4604 23520 4644
rect 24762 4632 24768 4684
rect 24820 4672 24826 4684
rect 24820 4644 25360 4672
rect 24820 4632 24826 4644
rect 23348 4576 23520 4604
rect 23348 4564 23354 4576
rect 23566 4564 23572 4616
rect 23624 4604 23630 4616
rect 23753 4607 23811 4613
rect 23753 4604 23765 4607
rect 23624 4576 23765 4604
rect 23624 4564 23630 4576
rect 23753 4573 23765 4576
rect 23799 4573 23811 4607
rect 23753 4567 23811 4573
rect 23842 4564 23848 4616
rect 23900 4604 23906 4616
rect 23900 4576 23945 4604
rect 23900 4564 23906 4576
rect 24486 4564 24492 4616
rect 24544 4604 24550 4616
rect 25332 4613 25360 4644
rect 26068 4613 26096 4780
rect 28166 4768 28172 4780
rect 28224 4768 28230 4820
rect 28258 4768 28264 4820
rect 28316 4808 28322 4820
rect 31386 4808 31392 4820
rect 28316 4780 31392 4808
rect 28316 4768 28322 4780
rect 31386 4768 31392 4780
rect 31444 4768 31450 4820
rect 34054 4768 34060 4820
rect 34112 4808 34118 4820
rect 38105 4811 38163 4817
rect 38105 4808 38117 4811
rect 34112 4780 38117 4808
rect 34112 4768 34118 4780
rect 38105 4777 38117 4780
rect 38151 4777 38163 4811
rect 38105 4771 38163 4777
rect 32306 4740 32312 4752
rect 28092 4712 32312 4740
rect 28092 4613 28120 4712
rect 32306 4700 32312 4712
rect 32364 4700 32370 4752
rect 31481 4675 31539 4681
rect 31481 4672 31493 4675
rect 31220 4644 31493 4672
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24544 4576 24685 4604
rect 24544 4564 24550 4576
rect 24673 4573 24685 4576
rect 24719 4604 24731 4607
rect 25225 4607 25283 4613
rect 25225 4604 25237 4607
rect 24719 4576 25237 4604
rect 24719 4573 24731 4576
rect 24673 4567 24731 4573
rect 25225 4573 25237 4576
rect 25271 4573 25283 4607
rect 25225 4567 25283 4573
rect 25317 4607 25375 4613
rect 25317 4573 25329 4607
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 26053 4607 26111 4613
rect 26053 4573 26065 4607
rect 26099 4604 26111 4607
rect 26329 4607 26387 4613
rect 26329 4604 26341 4607
rect 26099 4576 26341 4604
rect 26099 4573 26111 4576
rect 26053 4567 26111 4573
rect 26329 4573 26341 4576
rect 26375 4573 26387 4607
rect 26329 4567 26387 4573
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4573 28135 4607
rect 28077 4567 28135 4573
rect 30929 4607 30987 4613
rect 30929 4573 30941 4607
rect 30975 4600 30987 4607
rect 31220 4604 31248 4644
rect 31481 4641 31493 4644
rect 31527 4641 31539 4675
rect 31481 4635 31539 4641
rect 31386 4604 31392 4616
rect 31036 4600 31248 4604
rect 30975 4576 31248 4600
rect 31347 4576 31392 4604
rect 30975 4573 31064 4576
rect 30929 4572 31064 4573
rect 30929 4567 30987 4572
rect 31386 4564 31392 4576
rect 31444 4564 31450 4616
rect 38286 4604 38292 4616
rect 38247 4576 38292 4604
rect 38286 4564 38292 4576
rect 38344 4564 38350 4616
rect 20588 4508 20852 4536
rect 20588 4496 20594 4508
rect 21082 4496 21088 4548
rect 21140 4536 21146 4548
rect 22557 4539 22615 4545
rect 22557 4536 22569 4539
rect 21140 4508 22569 4536
rect 21140 4496 21146 4508
rect 22557 4505 22569 4508
rect 22603 4505 22615 4539
rect 22557 4499 22615 4505
rect 14918 4468 14924 4480
rect 8036 4440 14924 4468
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15930 4428 15936 4480
rect 15988 4468 15994 4480
rect 16025 4471 16083 4477
rect 16025 4468 16037 4471
rect 15988 4440 16037 4468
rect 15988 4428 15994 4440
rect 16025 4437 16037 4440
rect 16071 4437 16083 4471
rect 16025 4431 16083 4437
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 19886 4468 19892 4480
rect 17368 4440 19892 4468
rect 17368 4428 17374 4440
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 21358 4468 21364 4480
rect 20036 4440 21364 4468
rect 20036 4428 20042 4440
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 21634 4428 21640 4480
rect 21692 4468 21698 4480
rect 21913 4471 21971 4477
rect 21913 4468 21925 4471
rect 21692 4440 21925 4468
rect 21692 4428 21698 4440
rect 21913 4437 21925 4440
rect 21959 4437 21971 4471
rect 21913 4431 21971 4437
rect 22002 4428 22008 4480
rect 22060 4468 22066 4480
rect 23106 4468 23112 4480
rect 22060 4440 23112 4468
rect 22060 4428 22066 4440
rect 23106 4428 23112 4440
rect 23164 4428 23170 4480
rect 23584 4468 23612 4564
rect 23658 4496 23664 4548
rect 23716 4536 23722 4548
rect 25409 4539 25467 4545
rect 25409 4536 25421 4539
rect 23716 4508 25421 4536
rect 23716 4496 23722 4508
rect 25409 4505 25421 4508
rect 25455 4505 25467 4539
rect 25409 4499 25467 4505
rect 30760 4508 31754 4536
rect 24578 4468 24584 4480
rect 23584 4440 24584 4468
rect 24578 4428 24584 4440
rect 24636 4468 24642 4480
rect 24762 4468 24768 4480
rect 24636 4440 24768 4468
rect 24636 4428 24642 4440
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 25038 4468 25044 4480
rect 24999 4440 25044 4468
rect 25038 4428 25044 4440
rect 25096 4428 25102 4480
rect 30760 4477 30788 4508
rect 30745 4471 30803 4477
rect 30745 4437 30757 4471
rect 30791 4437 30803 4471
rect 31726 4468 31754 4508
rect 34422 4468 34428 4480
rect 31726 4440 34428 4468
rect 30745 4431 30803 4437
rect 34422 4428 34428 4440
rect 34480 4428 34486 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2038 4224 2044 4276
rect 2096 4264 2102 4276
rect 4890 4264 4896 4276
rect 2096 4236 4896 4264
rect 2096 4224 2102 4236
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 3160 4137 3188 4236
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5074 4224 5080 4276
rect 5132 4264 5138 4276
rect 12894 4264 12900 4276
rect 5132 4236 12900 4264
rect 5132 4224 5138 4236
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 16850 4264 16856 4276
rect 13872 4236 16856 4264
rect 13872 4224 13878 4236
rect 3418 4196 3424 4208
rect 3379 4168 3424 4196
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 6454 4196 6460 4208
rect 4646 4168 6460 4196
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6822 4196 6828 4208
rect 6656 4168 6828 4196
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 3145 4131 3203 4137
rect 2547 4100 2774 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 2746 4060 2774 4100
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5776 4100 5825 4128
rect 5776 4088 5782 4100
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6178 4128 6184 4140
rect 5951 4100 6184 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6656 4137 6684 4168
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 10870 4196 10876 4208
rect 6972 4168 7406 4196
rect 10810 4168 10876 4196
rect 6972 4156 6978 4168
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 13998 4196 14004 4208
rect 13202 4168 14004 4196
rect 13998 4156 14004 4168
rect 14056 4156 14062 4208
rect 14461 4199 14519 4205
rect 14461 4165 14473 4199
rect 14507 4196 14519 4199
rect 14568 4196 14596 4236
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 17236 4236 19380 4264
rect 17236 4196 17264 4236
rect 14507 4168 14596 4196
rect 15686 4168 17264 4196
rect 17313 4199 17371 4205
rect 14507 4165 14519 4168
rect 14461 4159 14519 4165
rect 17313 4165 17325 4199
rect 17359 4196 17371 4199
rect 19150 4196 19156 4208
rect 17359 4168 18092 4196
rect 17359 4165 17371 4168
rect 17313 4159 17371 4165
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8846 4128 8852 4140
rect 8352 4100 8852 4128
rect 8352 4088 8358 4100
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 14182 4128 14188 4140
rect 14143 4100 14188 4128
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 18064 4128 18092 4168
rect 19076 4168 19156 4196
rect 19076 4128 19104 4168
rect 19150 4156 19156 4168
rect 19208 4156 19214 4208
rect 19352 4196 19380 4236
rect 19426 4224 19432 4276
rect 19484 4264 19490 4276
rect 19889 4267 19947 4273
rect 19889 4264 19901 4267
rect 19484 4236 19901 4264
rect 19484 4224 19490 4236
rect 19889 4233 19901 4236
rect 19935 4233 19947 4267
rect 20346 4264 20352 4276
rect 20307 4236 20352 4264
rect 19889 4227 19947 4233
rect 20346 4224 20352 4236
rect 20404 4224 20410 4276
rect 20714 4224 20720 4276
rect 20772 4264 20778 4276
rect 21085 4267 21143 4273
rect 21085 4264 21097 4267
rect 20772 4236 21097 4264
rect 20772 4224 20778 4236
rect 21085 4233 21097 4236
rect 21131 4233 21143 4267
rect 22002 4264 22008 4276
rect 21085 4227 21143 4233
rect 21836 4236 22008 4264
rect 21836 4196 21864 4236
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 22738 4264 22744 4276
rect 22699 4236 22744 4264
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 23106 4224 23112 4276
rect 23164 4264 23170 4276
rect 25317 4267 25375 4273
rect 25317 4264 25329 4267
rect 23164 4236 25329 4264
rect 23164 4224 23170 4236
rect 25317 4233 25329 4236
rect 25363 4233 25375 4267
rect 25317 4227 25375 4233
rect 19352 4168 21864 4196
rect 21928 4168 22140 4196
rect 19978 4128 19984 4140
rect 18064 4100 19104 4128
rect 19168 4100 19984 4128
rect 4706 4060 4712 4072
rect 2746 4032 4712 4060
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4060 4951 4063
rect 5258 4060 5264 4072
rect 4939 4032 5264 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5994 4020 6000 4072
rect 6052 4060 6058 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6052 4032 6929 4060
rect 6052 4020 6058 4032
rect 1762 3992 1768 4004
rect 1723 3964 1768 3992
rect 1762 3952 1768 3964
rect 1820 3952 1826 4004
rect 6638 3992 6644 4004
rect 4816 3964 6644 3992
rect 2593 3927 2651 3933
rect 2593 3893 2605 3927
rect 2639 3924 2651 3927
rect 4816 3924 4844 3964
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 6748 3936 6776 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 9122 4060 9128 4072
rect 7708 4032 9128 4060
rect 7708 4020 7714 4032
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9674 4060 9680 4072
rect 9355 4032 9680 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9674 4020 9680 4032
rect 9732 4060 9738 4072
rect 10962 4060 10968 4072
rect 9732 4032 10968 4060
rect 9732 4020 9738 4032
rect 10962 4020 10968 4032
rect 11020 4060 11026 4072
rect 11698 4060 11704 4072
rect 11020 4032 11704 4060
rect 11020 4020 11026 4032
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11808 4032 11989 4060
rect 11057 3995 11115 4001
rect 11057 3961 11069 3995
rect 11103 3992 11115 3995
rect 11808 3992 11836 4032
rect 11977 4029 11989 4032
rect 12023 4060 12035 4063
rect 12023 4032 13124 4060
rect 12023 4029 12035 4032
rect 11977 4023 12035 4029
rect 11103 3964 11836 3992
rect 13096 3992 13124 4032
rect 13262 4020 13268 4072
rect 13320 4060 13326 4072
rect 13725 4063 13783 4069
rect 13725 4060 13737 4063
rect 13320 4032 13737 4060
rect 13320 4020 13326 4032
rect 13725 4029 13737 4032
rect 13771 4060 13783 4063
rect 14090 4060 14096 4072
rect 13771 4032 14096 4060
rect 13771 4029 13783 4032
rect 13725 4023 13783 4029
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 14550 4020 14556 4072
rect 14608 4060 14614 4072
rect 17221 4063 17279 4069
rect 14608 4032 15976 4060
rect 14608 4020 14614 4032
rect 13814 3992 13820 4004
rect 13096 3964 13820 3992
rect 11103 3961 11115 3964
rect 11057 3955 11115 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 2639 3896 4844 3924
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 6730 3884 6736 3936
rect 6788 3884 6794 3936
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 9398 3924 9404 3936
rect 8435 3896 9404 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9572 3927 9630 3933
rect 9572 3893 9584 3927
rect 9618 3924 9630 3927
rect 11606 3924 11612 3936
rect 9618 3896 11612 3924
rect 9618 3893 9630 3896
rect 9572 3887 9630 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12434 3924 12440 3936
rect 12032 3896 12440 3924
rect 12032 3884 12038 3896
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 15948 3933 15976 4032
rect 17221 4029 17233 4063
rect 17267 4060 17279 4063
rect 17586 4060 17592 4072
rect 17267 4032 17592 4060
rect 17267 4029 17279 4032
rect 17221 4023 17279 4029
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 17678 4020 17684 4072
rect 17736 4060 17742 4072
rect 18233 4063 18291 4069
rect 18233 4060 18245 4063
rect 17736 4032 18245 4060
rect 17736 4020 17742 4032
rect 18233 4029 18245 4032
rect 18279 4060 18291 4063
rect 19058 4060 19064 4072
rect 18279 4032 19064 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 16758 3952 16764 4004
rect 16816 3992 16822 4004
rect 19168 3992 19196 4100
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4128 21051 4131
rect 21928 4128 21956 4168
rect 21039 4100 21956 4128
rect 22005 4131 22063 4137
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 19429 4063 19487 4069
rect 19429 4029 19441 4063
rect 19475 4060 19487 4063
rect 21174 4060 21180 4072
rect 19475 4032 21180 4060
rect 19475 4029 19487 4032
rect 19429 4023 19487 4029
rect 16816 3964 19196 3992
rect 19260 3992 19288 4023
rect 21174 4020 21180 4032
rect 21232 4020 21238 4072
rect 21266 4020 21272 4072
rect 21324 4060 21330 4072
rect 22020 4060 22048 4091
rect 21324 4032 22048 4060
rect 22112 4060 22140 4168
rect 23676 4168 24716 4196
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 22649 4131 22707 4137
rect 22649 4128 22661 4131
rect 22244 4100 22661 4128
rect 22244 4088 22250 4100
rect 22649 4097 22661 4100
rect 22695 4128 22707 4131
rect 23293 4131 23351 4137
rect 23293 4128 23305 4131
rect 22695 4100 23305 4128
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 23293 4097 23305 4100
rect 23339 4128 23351 4131
rect 23676 4128 23704 4168
rect 23339 4100 23704 4128
rect 23339 4097 23351 4100
rect 23293 4091 23351 4097
rect 23750 4088 23756 4140
rect 23808 4128 23814 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 23808 4100 23949 4128
rect 23808 4088 23814 4100
rect 23937 4097 23949 4100
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4097 24639 4131
rect 24688 4128 24716 4168
rect 37182 4156 37188 4208
rect 37240 4196 37246 4208
rect 38105 4199 38163 4205
rect 38105 4196 38117 4199
rect 37240 4168 38117 4196
rect 37240 4156 37246 4168
rect 38105 4165 38117 4168
rect 38151 4165 38163 4199
rect 38105 4159 38163 4165
rect 25225 4131 25283 4137
rect 25225 4128 25237 4131
rect 24688 4100 25237 4128
rect 24581 4091 24639 4097
rect 25225 4097 25237 4100
rect 25271 4128 25283 4131
rect 25774 4128 25780 4140
rect 25271 4100 25780 4128
rect 25271 4097 25283 4100
rect 25225 4091 25283 4097
rect 23014 4060 23020 4072
rect 22112 4032 23020 4060
rect 21324 4020 21330 4032
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 23198 4020 23204 4072
rect 23256 4060 23262 4072
rect 24596 4060 24624 4091
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 27338 4128 27344 4140
rect 27299 4100 27344 4128
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 25130 4060 25136 4072
rect 23256 4032 25136 4060
rect 23256 4020 23262 4032
rect 25130 4020 25136 4032
rect 25188 4020 25194 4072
rect 20806 3992 20812 4004
rect 19260 3964 20812 3992
rect 16816 3952 16822 3964
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 21726 3952 21732 4004
rect 21784 3992 21790 4004
rect 22097 3995 22155 4001
rect 22097 3992 22109 3995
rect 21784 3964 22109 3992
rect 21784 3952 21790 3964
rect 22097 3961 22109 3964
rect 22143 3961 22155 3995
rect 22097 3955 22155 3961
rect 24762 3952 24768 4004
rect 24820 3992 24826 4004
rect 26053 3995 26111 4001
rect 26053 3992 26065 3995
rect 24820 3964 26065 3992
rect 24820 3952 24826 3964
rect 26053 3961 26065 3964
rect 26099 3961 26111 3995
rect 26053 3955 26111 3961
rect 26878 3952 26884 4004
rect 26936 3992 26942 4004
rect 26936 3964 35894 3992
rect 26936 3952 26942 3964
rect 15933 3927 15991 3933
rect 15933 3893 15945 3927
rect 15979 3924 15991 3927
rect 16298 3924 16304 3936
rect 15979 3896 16304 3924
rect 15979 3893 15991 3896
rect 15933 3887 15991 3893
rect 16298 3884 16304 3896
rect 16356 3924 16362 3936
rect 21634 3924 21640 3936
rect 16356 3896 21640 3924
rect 16356 3884 16362 3896
rect 21634 3884 21640 3896
rect 21692 3884 21698 3936
rect 23382 3924 23388 3936
rect 23343 3896 23388 3924
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 24026 3924 24032 3936
rect 23987 3896 24032 3924
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24118 3884 24124 3936
rect 24176 3924 24182 3936
rect 24673 3927 24731 3933
rect 24673 3924 24685 3927
rect 24176 3896 24685 3924
rect 24176 3884 24182 3896
rect 24673 3893 24685 3896
rect 24719 3893 24731 3927
rect 24673 3887 24731 3893
rect 26694 3884 26700 3936
rect 26752 3924 26758 3936
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 26752 3896 27169 3924
rect 26752 3884 26758 3896
rect 27157 3893 27169 3896
rect 27203 3893 27215 3927
rect 35866 3924 35894 3964
rect 38197 3927 38255 3933
rect 38197 3924 38209 3927
rect 35866 3896 38209 3924
rect 27157 3887 27215 3893
rect 38197 3893 38209 3896
rect 38243 3893 38255 3927
rect 38197 3887 38255 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 2498 3720 2504 3732
rect 2271 3692 2504 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2240 3516 2268 3683
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 6086 3720 6092 3732
rect 4120 3692 6092 3720
rect 4120 3680 4126 3692
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 9769 3723 9827 3729
rect 9769 3689 9781 3723
rect 9815 3720 9827 3723
rect 9858 3720 9864 3732
rect 9815 3692 9864 3720
rect 9815 3689 9827 3692
rect 9769 3683 9827 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10584 3723 10642 3729
rect 10584 3689 10596 3723
rect 10630 3720 10642 3723
rect 11974 3720 11980 3732
rect 10630 3692 11980 3720
rect 10630 3689 10642 3692
rect 10584 3683 10642 3689
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12308 3692 13001 3720
rect 12308 3680 12314 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 12989 3683 13047 3689
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13228 3692 13645 3720
rect 13228 3680 13234 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13633 3683 13691 3689
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 19886 3720 19892 3732
rect 14608 3692 19892 3720
rect 14608 3680 14614 3692
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 20162 3720 20168 3732
rect 20123 3692 20168 3720
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 24670 3720 24676 3732
rect 20680 3692 24676 3720
rect 20680 3680 20686 3692
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 25866 3680 25872 3732
rect 25924 3720 25930 3732
rect 25961 3723 26019 3729
rect 25961 3720 25973 3723
rect 25924 3692 25973 3720
rect 25924 3680 25930 3692
rect 25961 3689 25973 3692
rect 26007 3689 26019 3723
rect 37734 3720 37740 3732
rect 25961 3683 26019 3689
rect 28966 3692 37740 3720
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3652 3387 3655
rect 4338 3652 4344 3664
rect 3375 3624 4344 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 4338 3612 4344 3624
rect 4396 3612 4402 3664
rect 7006 3652 7012 3664
rect 6380 3624 7012 3652
rect 6380 3584 6408 3624
rect 7006 3612 7012 3624
rect 7064 3612 7070 3664
rect 7193 3655 7251 3661
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 8570 3652 8576 3664
rect 7239 3624 8576 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 8570 3612 8576 3624
rect 8628 3612 8634 3664
rect 11606 3612 11612 3664
rect 11664 3652 11670 3664
rect 13538 3652 13544 3664
rect 11664 3624 13544 3652
rect 11664 3612 11670 3624
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 14274 3612 14280 3664
rect 14332 3652 14338 3664
rect 18966 3652 18972 3664
rect 14332 3624 18972 3652
rect 14332 3612 14338 3624
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 20070 3652 20076 3664
rect 19076 3624 20076 3652
rect 4448 3556 6408 3584
rect 1627 3488 2268 3516
rect 2593 3519 2651 3525
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 4338 3516 4344 3528
rect 3283 3488 4344 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 2608 3448 2636 3479
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4448 3448 4476 3556
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 10321 3587 10379 3593
rect 6788 3556 9720 3584
rect 6788 3544 6794 3556
rect 4525 3519 4583 3525
rect 4525 3485 4537 3519
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6822 3516 6828 3528
rect 6595 3488 6828 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 2608 3420 4476 3448
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3380 2743 3383
rect 4430 3380 4436 3392
rect 2731 3352 4436 3380
rect 2731 3349 2743 3352
rect 2685 3343 2743 3349
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4547 3380 4575 3479
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7650 3516 7656 3528
rect 7147 3488 7656 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 8294 3516 8300 3528
rect 7791 3488 8300 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 9582 3516 9588 3528
rect 8435 3488 9588 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9692 3525 9720 3556
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 11790 3584 11796 3596
rect 10367 3556 11796 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 12342 3584 12348 3596
rect 12303 3556 12348 3584
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 15657 3587 15715 3593
rect 15657 3553 15669 3587
rect 15703 3584 15715 3587
rect 16114 3584 16120 3596
rect 15703 3556 16120 3584
rect 15703 3553 15715 3556
rect 15657 3547 15715 3553
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 19076 3584 19104 3624
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 20346 3612 20352 3664
rect 20404 3652 20410 3664
rect 21453 3655 21511 3661
rect 21453 3652 21465 3655
rect 20404 3624 21465 3652
rect 20404 3612 20410 3624
rect 21453 3621 21465 3624
rect 21499 3621 21511 3655
rect 22094 3652 22100 3664
rect 22055 3624 22100 3652
rect 21453 3615 21511 3621
rect 22094 3612 22100 3624
rect 22152 3612 22158 3664
rect 28966 3652 28994 3692
rect 37734 3680 37740 3692
rect 37792 3680 37798 3732
rect 37553 3655 37611 3661
rect 37553 3652 37565 3655
rect 22204 3624 28994 3652
rect 35866 3624 37565 3652
rect 17000 3556 19104 3584
rect 17000 3544 17006 3556
rect 19334 3544 19340 3596
rect 19392 3584 19398 3596
rect 19521 3587 19579 3593
rect 19521 3584 19533 3587
rect 19392 3556 19533 3584
rect 19392 3544 19398 3556
rect 19521 3553 19533 3556
rect 19567 3553 19579 3587
rect 19521 3547 19579 3553
rect 20530 3544 20536 3596
rect 20588 3544 20594 3596
rect 20806 3584 20812 3596
rect 20767 3556 20812 3584
rect 20806 3544 20812 3556
rect 20864 3544 20870 3596
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 22204 3584 22232 3624
rect 25038 3584 25044 3596
rect 21968 3556 22232 3584
rect 22388 3556 25044 3584
rect 21968 3544 21974 3556
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12897 3519 12955 3525
rect 12897 3516 12909 3519
rect 12032 3488 12909 3516
rect 12032 3476 12038 3488
rect 12897 3485 12909 3488
rect 12943 3516 12955 3519
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 12943 3488 13553 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 16758 3516 16764 3528
rect 16719 3488 16764 3516
rect 13541 3479 13599 3485
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3516 16911 3519
rect 17034 3516 17040 3528
rect 16899 3488 17040 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18690 3516 18696 3528
rect 18463 3488 18696 3516
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20548 3516 20576 3544
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 20119 3488 20484 3516
rect 20548 3488 20729 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 4798 3408 4804 3460
rect 4856 3448 4862 3460
rect 4856 3420 4901 3448
rect 6026 3420 6224 3448
rect 4856 3408 4862 3420
rect 4890 3380 4896 3392
rect 4547 3352 4896 3380
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 6196 3380 6224 3420
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 6696 3420 11086 3448
rect 6696 3408 6702 3420
rect 12158 3408 12164 3460
rect 12216 3448 12222 3460
rect 14274 3448 14280 3460
rect 12216 3420 14280 3448
rect 12216 3408 12222 3420
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 14461 3451 14519 3457
rect 14461 3417 14473 3451
rect 14507 3417 14519 3451
rect 14461 3411 14519 3417
rect 7006 3380 7012 3392
rect 6196 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7837 3383 7895 3389
rect 7837 3349 7849 3383
rect 7883 3380 7895 3383
rect 8662 3380 8668 3392
rect 7883 3352 8668 3380
rect 7883 3349 7895 3352
rect 7837 3343 7895 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 13354 3380 13360 3392
rect 11296 3352 13360 3380
rect 11296 3340 11302 3352
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 14476 3380 14504 3411
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 15105 3451 15163 3457
rect 14608 3420 14653 3448
rect 14608 3408 14614 3420
rect 15105 3417 15117 3451
rect 15151 3448 15163 3451
rect 15194 3448 15200 3460
rect 15151 3420 15200 3448
rect 15151 3417 15163 3420
rect 15105 3411 15163 3417
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 15749 3451 15807 3457
rect 15749 3417 15761 3451
rect 15795 3417 15807 3451
rect 15749 3411 15807 3417
rect 14734 3380 14740 3392
rect 14476 3352 14740 3380
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 15764 3380 15792 3411
rect 15838 3408 15844 3460
rect 15896 3448 15902 3460
rect 16301 3451 16359 3457
rect 16301 3448 16313 3451
rect 15896 3420 16313 3448
rect 15896 3408 15902 3420
rect 16301 3417 16313 3420
rect 16347 3417 16359 3451
rect 17770 3448 17776 3460
rect 17731 3420 17776 3448
rect 16301 3411 16359 3417
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 17865 3451 17923 3457
rect 17865 3417 17877 3451
rect 17911 3417 17923 3451
rect 18708 3448 18736 3476
rect 19702 3448 19708 3460
rect 18708 3420 19708 3448
rect 17865 3411 17923 3417
rect 17678 3380 17684 3392
rect 15764 3352 17684 3380
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 17880 3380 17908 3411
rect 19702 3408 19708 3420
rect 19760 3408 19766 3460
rect 20070 3380 20076 3392
rect 17880 3352 20076 3380
rect 20070 3340 20076 3352
rect 20128 3340 20134 3392
rect 20456 3380 20484 3488
rect 20717 3485 20729 3488
rect 20763 3485 20775 3519
rect 21358 3516 21364 3528
rect 21319 3488 21364 3516
rect 20717 3479 20775 3485
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 22005 3519 22063 3525
rect 22005 3516 22017 3519
rect 21508 3488 22017 3516
rect 21508 3476 21514 3488
rect 22005 3485 22017 3488
rect 22051 3485 22063 3519
rect 22005 3479 22063 3485
rect 20530 3408 20536 3460
rect 20588 3448 20594 3460
rect 21082 3448 21088 3460
rect 20588 3420 21088 3448
rect 20588 3408 20594 3420
rect 21082 3408 21088 3420
rect 21140 3408 21146 3460
rect 22388 3448 22416 3556
rect 25038 3544 25044 3556
rect 25096 3544 25102 3596
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 22520 3488 22661 3516
rect 22520 3476 22526 3488
rect 22649 3485 22661 3488
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 22741 3519 22799 3525
rect 22741 3485 22753 3519
rect 22787 3516 22799 3519
rect 23477 3519 23535 3525
rect 22787 3488 23428 3516
rect 22787 3485 22799 3488
rect 22741 3479 22799 3485
rect 21192 3420 22416 3448
rect 23400 3448 23428 3488
rect 23477 3485 23489 3519
rect 23523 3516 23535 3519
rect 24210 3516 24216 3528
rect 23523 3488 24216 3516
rect 23523 3485 23535 3488
rect 23477 3479 23535 3485
rect 24210 3476 24216 3488
rect 24268 3476 24274 3528
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 25130 3476 25136 3528
rect 25188 3516 25194 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 25188 3488 25237 3516
rect 25188 3476 25194 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25774 3476 25780 3528
rect 25832 3516 25838 3528
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 25832 3488 25881 3516
rect 25832 3476 25838 3488
rect 25869 3485 25881 3488
rect 25915 3516 25927 3519
rect 26513 3519 26571 3525
rect 26513 3516 26525 3519
rect 25915 3488 26525 3516
rect 25915 3485 25927 3488
rect 25869 3479 25927 3485
rect 26513 3485 26525 3488
rect 26559 3485 26571 3519
rect 26513 3479 26571 3485
rect 27341 3519 27399 3525
rect 27341 3485 27353 3519
rect 27387 3485 27399 3519
rect 27982 3516 27988 3528
rect 27943 3488 27988 3516
rect 27341 3479 27399 3485
rect 27356 3448 27384 3479
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 23400 3420 27384 3448
rect 21192 3380 21220 3420
rect 27430 3408 27436 3460
rect 27488 3448 27494 3460
rect 35866 3448 35894 3624
rect 37553 3621 37565 3624
rect 37599 3621 37611 3655
rect 37553 3615 37611 3621
rect 37918 3476 37924 3528
rect 37976 3516 37982 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37976 3488 38025 3516
rect 37976 3476 37982 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 27488 3420 35894 3448
rect 37369 3451 37427 3457
rect 27488 3408 27494 3420
rect 37369 3417 37381 3451
rect 37415 3448 37427 3451
rect 37415 3420 38056 3448
rect 37415 3417 37427 3420
rect 37369 3411 37427 3417
rect 38028 3392 38056 3420
rect 20456 3352 21220 3380
rect 22186 3340 22192 3392
rect 22244 3380 22250 3392
rect 23293 3383 23351 3389
rect 23293 3380 23305 3383
rect 22244 3352 23305 3380
rect 22244 3340 22250 3352
rect 23293 3349 23305 3352
rect 23339 3349 23351 3383
rect 23293 3343 23351 3349
rect 23474 3340 23480 3392
rect 23532 3380 23538 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 23532 3352 24685 3380
rect 23532 3340 23538 3352
rect 24673 3349 24685 3352
rect 24719 3349 24731 3383
rect 24673 3343 24731 3349
rect 24854 3340 24860 3392
rect 24912 3380 24918 3392
rect 25317 3383 25375 3389
rect 25317 3380 25329 3383
rect 24912 3352 25329 3380
rect 24912 3340 24918 3352
rect 25317 3349 25329 3352
rect 25363 3349 25375 3383
rect 26602 3380 26608 3392
rect 26563 3352 26608 3380
rect 25317 3343 25375 3349
rect 26602 3340 26608 3352
rect 26660 3340 26666 3392
rect 27154 3380 27160 3392
rect 27115 3352 27160 3380
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 27798 3380 27804 3392
rect 27759 3352 27804 3380
rect 27798 3340 27804 3352
rect 27856 3340 27862 3392
rect 38010 3340 38016 3392
rect 38068 3340 38074 3392
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3329 3179 3387 3185
rect 3329 3145 3341 3179
rect 3375 3176 3387 3179
rect 4430 3176 4436 3188
rect 3375 3148 4436 3176
rect 3375 3145 3387 3148
rect 3329 3139 3387 3145
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 5442 3176 5448 3188
rect 5307 3148 5448 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6825 3179 6883 3185
rect 6825 3145 6837 3179
rect 6871 3176 6883 3179
rect 7558 3176 7564 3188
rect 6871 3148 7564 3176
rect 6871 3145 6883 3148
rect 6825 3139 6883 3145
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8168 3148 8769 3176
rect 8168 3136 8174 3148
rect 8757 3145 8769 3148
rect 8803 3145 8815 3179
rect 10410 3176 10416 3188
rect 10371 3148 10416 3176
rect 8757 3139 8815 3145
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 11057 3179 11115 3185
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 12802 3176 12808 3188
rect 11103 3148 12808 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 14737 3179 14795 3185
rect 13504 3148 14688 3176
rect 13504 3136 13510 3148
rect 2406 3108 2412 3120
rect 1596 3080 2412 3108
rect 1596 3049 1624 3080
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 4617 3111 4675 3117
rect 3252 3080 4568 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 1581 3003 1639 3009
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 3252 3049 3280 3080
rect 4540 3049 4568 3080
rect 4617 3077 4629 3111
rect 4663 3108 4675 3111
rect 5534 3108 5540 3120
rect 4663 3080 5540 3108
rect 4663 3077 4675 3080
rect 4617 3071 4675 3077
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 5905 3111 5963 3117
rect 5905 3077 5917 3111
rect 5951 3108 5963 3111
rect 6638 3108 6644 3120
rect 5951 3080 6644 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 7248 3080 12558 3108
rect 13924 3080 14596 3108
rect 7248 3068 7254 3080
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 5166 3040 5172 3052
rect 4571 3012 5172 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 14 2864 20 2916
rect 72 2904 78 2916
rect 2501 2907 2559 2913
rect 2501 2904 2513 2907
rect 72 2876 2513 2904
rect 72 2864 78 2876
rect 2501 2873 2513 2876
rect 2547 2873 2559 2907
rect 2501 2867 2559 2873
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 716 2808 1777 2836
rect 716 2796 722 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 3896 2836 3924 3003
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 5868 3012 5913 3040
rect 5868 3000 5874 3012
rect 6546 3000 6552 3052
rect 6604 3040 6610 3052
rect 6741 3049 6799 3055
rect 6604 3038 6684 3040
rect 6741 3038 6753 3049
rect 6604 3015 6753 3038
rect 6787 3015 6799 3049
rect 7374 3040 7380 3052
rect 6604 3012 6799 3015
rect 7287 3012 7380 3040
rect 6604 3000 6610 3012
rect 6656 3010 6799 3012
rect 6741 3009 6799 3010
rect 7374 3000 7380 3012
rect 7432 3040 7438 3052
rect 7432 3012 7604 3040
rect 7432 3000 7438 3012
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 5626 2972 5632 2984
rect 4019 2944 5632 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 6512 2944 7481 2972
rect 6512 2932 6518 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 4430 2864 4436 2916
rect 4488 2904 4494 2916
rect 7190 2904 7196 2916
rect 4488 2876 7196 2904
rect 4488 2864 4494 2876
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 7576 2904 7604 3012
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7892 3012 8033 3040
rect 7892 3000 7898 3012
rect 8021 3009 8033 3012
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8260 3012 8677 3040
rect 8260 3000 8266 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 9324 2972 9352 3003
rect 10226 3000 10232 3052
rect 10284 3040 10290 3052
rect 10321 3043 10379 3049
rect 10321 3040 10333 3043
rect 10284 3012 10333 3040
rect 10284 3000 10290 3012
rect 10321 3009 10333 3012
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10744 3012 10977 3040
rect 10744 3000 10750 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 11790 3040 11796 3052
rect 11751 3012 11796 3040
rect 10965 3003 11023 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 7984 2944 9352 2972
rect 7984 2932 7990 2944
rect 9324 2904 9352 2944
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 11054 2972 11060 2984
rect 9447 2944 11060 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11480 2944 12081 2972
rect 11480 2932 11486 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 13538 2972 13544 2984
rect 13451 2944 13544 2972
rect 12069 2935 12127 2941
rect 13538 2932 13544 2944
rect 13596 2972 13602 2984
rect 13722 2972 13728 2984
rect 13596 2944 13728 2972
rect 13596 2932 13602 2944
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 11238 2904 11244 2916
rect 7576 2876 8248 2904
rect 9324 2876 11244 2904
rect 5718 2836 5724 2848
rect 3896 2808 5724 2836
rect 1765 2799 1823 2805
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 6420 2808 8125 2836
rect 6420 2796 6426 2808
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 8220 2836 8248 2876
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 12710 2836 12716 2848
rect 8220 2808 12716 2836
rect 8113 2799 8171 2805
rect 12710 2796 12716 2808
rect 12768 2836 12774 2848
rect 13924 2836 13952 3080
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14016 2904 14044 3003
rect 14568 2972 14596 3080
rect 14660 3049 14688 3148
rect 14737 3145 14749 3179
rect 14783 3176 14795 3179
rect 15102 3176 15108 3188
rect 14783 3148 15108 3176
rect 14783 3145 14795 3148
rect 14737 3139 14795 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 16022 3176 16028 3188
rect 15983 3148 16028 3176
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 16390 3136 16396 3188
rect 16448 3176 16454 3188
rect 18414 3176 18420 3188
rect 16448 3148 17264 3176
rect 18375 3148 18420 3176
rect 16448 3136 16454 3148
rect 14918 3068 14924 3120
rect 14976 3108 14982 3120
rect 16482 3108 16488 3120
rect 14976 3080 16488 3108
rect 14976 3068 14982 3080
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 15297 3043 15355 3049
rect 15297 3009 15309 3043
rect 15343 3040 15355 3043
rect 15396 3040 15424 3080
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 17236 3117 17264 3148
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 18506 3136 18512 3188
rect 18564 3176 18570 3188
rect 19061 3179 19119 3185
rect 19061 3176 19073 3179
rect 18564 3148 19073 3176
rect 18564 3136 18570 3148
rect 19061 3145 19073 3148
rect 19107 3145 19119 3179
rect 19061 3139 19119 3145
rect 19150 3136 19156 3188
rect 19208 3176 19214 3188
rect 19705 3179 19763 3185
rect 19705 3176 19717 3179
rect 19208 3148 19717 3176
rect 19208 3136 19214 3148
rect 19705 3145 19717 3148
rect 19751 3145 19763 3179
rect 20806 3176 20812 3188
rect 19705 3139 19763 3145
rect 20081 3148 20812 3176
rect 17221 3111 17279 3117
rect 17221 3077 17233 3111
rect 17267 3077 17279 3111
rect 17221 3071 17279 3077
rect 17313 3111 17371 3117
rect 17313 3077 17325 3111
rect 17359 3108 17371 3111
rect 20081 3108 20109 3148
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 27801 3179 27859 3185
rect 27801 3176 27813 3179
rect 21416 3148 27813 3176
rect 21416 3136 21422 3148
rect 27801 3145 27813 3148
rect 27847 3145 27859 3179
rect 27801 3139 27859 3145
rect 30742 3136 30748 3188
rect 30800 3176 30806 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 30800 3148 36737 3176
rect 30800 3136 30806 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 22370 3108 22376 3120
rect 17359 3080 20109 3108
rect 22066 3080 22376 3108
rect 17359 3077 17371 3080
rect 17313 3071 17371 3077
rect 15343 3012 15424 3040
rect 15933 3043 15991 3049
rect 15343 3009 15355 3012
rect 15297 3003 15355 3009
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16758 3040 16764 3052
rect 15979 3012 16764 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 15948 2972 15976 3003
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 18322 3040 18328 3052
rect 18283 3012 18328 3040
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 18966 3040 18972 3052
rect 18927 3012 18972 3040
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 19610 3000 19616 3052
rect 19668 3047 19674 3052
rect 19668 3038 19679 3047
rect 19668 3010 19711 3038
rect 19668 3001 19679 3010
rect 19668 3000 19674 3001
rect 20162 3000 20168 3052
rect 20220 3038 20226 3052
rect 20257 3043 20315 3049
rect 20257 3038 20269 3043
rect 20220 3010 20269 3038
rect 20220 3000 20226 3010
rect 20257 3009 20269 3010
rect 20303 3009 20315 3043
rect 20257 3003 20315 3009
rect 20346 3000 20352 3052
rect 20404 3040 20410 3052
rect 21085 3043 21143 3049
rect 20404 3012 20449 3040
rect 20404 3000 20410 3012
rect 21085 3009 21097 3043
rect 21131 3040 21143 3043
rect 22066 3040 22094 3080
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 24670 3068 24676 3120
rect 24728 3108 24734 3120
rect 24857 3111 24915 3117
rect 24857 3108 24869 3111
rect 24728 3080 24869 3108
rect 24728 3068 24734 3080
rect 24857 3077 24869 3080
rect 24903 3077 24915 3111
rect 25498 3108 25504 3120
rect 25459 3080 25504 3108
rect 24857 3071 24915 3077
rect 25498 3068 25504 3080
rect 25556 3068 25562 3120
rect 21131 3012 22094 3040
rect 22189 3043 22247 3049
rect 21131 3009 21143 3012
rect 21085 3003 21143 3009
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22646 3040 22652 3052
rect 22607 3012 22652 3040
rect 22189 3003 22247 3009
rect 14568 2944 15976 2972
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2972 17923 2975
rect 18230 2972 18236 2984
rect 17911 2944 18236 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 22204 2972 22232 3003
rect 22646 3000 22652 3012
rect 22704 3000 22710 3052
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 23937 3043 23995 3049
rect 23937 3009 23949 3043
rect 23983 3040 23995 3043
rect 24765 3043 24823 3049
rect 23983 3012 24164 3040
rect 23983 3009 23995 3012
rect 23937 3003 23995 3009
rect 19392 2944 22232 2972
rect 19392 2932 19398 2944
rect 22278 2932 22284 2984
rect 22336 2972 22342 2984
rect 22922 2972 22928 2984
rect 22336 2944 22928 2972
rect 22336 2932 22342 2944
rect 22922 2932 22928 2944
rect 22980 2932 22986 2984
rect 23492 2972 23520 3003
rect 24029 2975 24087 2981
rect 24029 2972 24041 2975
rect 23492 2944 24041 2972
rect 24029 2941 24041 2944
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 14016 2876 16712 2904
rect 12768 2808 13952 2836
rect 14093 2839 14151 2845
rect 12768 2796 12774 2808
rect 14093 2805 14105 2839
rect 14139 2836 14151 2839
rect 15286 2836 15292 2848
rect 14139 2808 15292 2836
rect 14139 2805 14151 2808
rect 14093 2799 14151 2805
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 16114 2836 16120 2848
rect 15712 2808 16120 2836
rect 15712 2796 15718 2808
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 16684 2836 16712 2876
rect 17310 2864 17316 2916
rect 17368 2904 17374 2916
rect 20530 2904 20536 2916
rect 17368 2876 20536 2904
rect 17368 2864 17374 2876
rect 20530 2864 20536 2876
rect 20588 2864 20594 2916
rect 22005 2907 22063 2913
rect 22005 2904 22017 2907
rect 20640 2876 22017 2904
rect 20640 2836 20668 2876
rect 22005 2873 22017 2876
rect 22051 2873 22063 2907
rect 24136 2904 24164 3012
rect 24765 3009 24777 3043
rect 24811 3040 24823 3043
rect 25314 3040 25320 3052
rect 24811 3012 25320 3040
rect 24811 3009 24823 3012
rect 24765 3003 24823 3009
rect 25314 3000 25320 3012
rect 25372 3000 25378 3052
rect 25406 3000 25412 3052
rect 25464 3040 25470 3052
rect 25464 3012 25509 3040
rect 25464 3000 25470 3012
rect 25682 3000 25688 3052
rect 25740 3040 25746 3052
rect 26237 3043 26295 3049
rect 26237 3040 26249 3043
rect 25740 3012 26249 3040
rect 25740 3000 25746 3012
rect 26237 3009 26249 3012
rect 26283 3009 26295 3043
rect 26237 3003 26295 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3040 27215 3043
rect 27982 3040 27988 3052
rect 27203 3012 27568 3040
rect 27943 3012 27988 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 24210 2932 24216 2984
rect 24268 2972 24274 2984
rect 27430 2972 27436 2984
rect 24268 2944 27436 2972
rect 24268 2932 24274 2944
rect 27430 2932 27436 2944
rect 27488 2932 27494 2984
rect 22005 2867 22063 2873
rect 22572 2876 24164 2904
rect 16684 2808 20668 2836
rect 20901 2839 20959 2845
rect 20901 2805 20913 2839
rect 20947 2836 20959 2839
rect 21818 2836 21824 2848
rect 20947 2808 21824 2836
rect 20947 2805 20959 2808
rect 20901 2799 20959 2805
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 21910 2796 21916 2848
rect 21968 2836 21974 2848
rect 22572 2836 22600 2876
rect 24578 2864 24584 2916
rect 24636 2904 24642 2916
rect 27540 2904 27568 3012
rect 27982 3000 27988 3012
rect 28040 3000 28046 3052
rect 36909 3043 36967 3049
rect 36909 3009 36921 3043
rect 36955 3040 36967 3043
rect 37734 3040 37740 3052
rect 36955 3012 37596 3040
rect 37695 3012 37740 3040
rect 36955 3009 36967 3012
rect 36909 3003 36967 3009
rect 37458 2972 37464 2984
rect 37419 2944 37464 2972
rect 37458 2932 37464 2944
rect 37516 2932 37522 2984
rect 37568 2972 37596 3012
rect 37734 3000 37740 3012
rect 37792 3000 37798 3052
rect 39298 2972 39304 2984
rect 37568 2944 39304 2972
rect 39298 2932 39304 2944
rect 39356 2932 39362 2984
rect 24636 2876 27568 2904
rect 24636 2864 24642 2876
rect 22738 2836 22744 2848
rect 21968 2808 22600 2836
rect 22699 2808 22744 2836
rect 21968 2796 21974 2808
rect 22738 2796 22744 2808
rect 22796 2796 22802 2848
rect 23290 2836 23296 2848
rect 23251 2808 23296 2836
rect 23290 2796 23296 2808
rect 23348 2796 23354 2848
rect 26050 2836 26056 2848
rect 26011 2808 26056 2836
rect 26050 2796 26056 2808
rect 26108 2796 26114 2848
rect 27246 2836 27252 2848
rect 27207 2808 27252 2836
rect 27246 2796 27252 2808
rect 27304 2796 27310 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7064 2604 7849 2632
rect 7064 2592 7070 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 9950 2632 9956 2644
rect 7837 2595 7895 2601
rect 8220 2604 9956 2632
rect 5442 2564 5448 2576
rect 2056 2536 5448 2564
rect 2056 2437 2084 2536
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 8220 2496 8248 2604
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 10505 2635 10563 2641
rect 10505 2632 10517 2635
rect 10192 2604 10517 2632
rect 10192 2592 10198 2604
rect 10505 2601 10517 2604
rect 10551 2601 10563 2635
rect 10505 2595 10563 2601
rect 12618 2592 12624 2644
rect 12676 2632 12682 2644
rect 13722 2632 13728 2644
rect 12676 2604 13728 2632
rect 12676 2592 12682 2604
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 14826 2632 14832 2644
rect 14787 2604 14832 2632
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 16114 2632 16120 2644
rect 16075 2604 16120 2632
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 16945 2635 17003 2641
rect 16945 2632 16957 2635
rect 16540 2604 16957 2632
rect 16540 2592 16546 2604
rect 16945 2601 16957 2604
rect 16991 2601 17003 2635
rect 16945 2595 17003 2601
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 17589 2635 17647 2641
rect 17589 2632 17601 2635
rect 17552 2604 17601 2632
rect 17552 2592 17558 2604
rect 17589 2601 17601 2604
rect 17635 2601 17647 2635
rect 17589 2595 17647 2601
rect 20165 2635 20223 2641
rect 20165 2601 20177 2635
rect 20211 2632 20223 2635
rect 20346 2632 20352 2644
rect 20211 2604 20352 2632
rect 20211 2601 20223 2604
rect 20165 2595 20223 2601
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 22646 2632 22652 2644
rect 22051 2604 22652 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 24302 2592 24308 2644
rect 24360 2632 24366 2644
rect 24581 2635 24639 2641
rect 24581 2632 24593 2635
rect 24360 2604 24593 2632
rect 24360 2592 24366 2604
rect 24581 2601 24593 2604
rect 24627 2601 24639 2635
rect 24581 2595 24639 2601
rect 25314 2592 25320 2644
rect 25372 2632 25378 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 25372 2604 27169 2632
rect 25372 2592 25378 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 28442 2632 28448 2644
rect 28403 2604 28448 2632
rect 27157 2595 27215 2601
rect 28442 2592 28448 2604
rect 28500 2592 28506 2644
rect 30466 2632 30472 2644
rect 30427 2604 30472 2632
rect 30466 2592 30472 2604
rect 30524 2592 30530 2644
rect 32306 2632 32312 2644
rect 32267 2604 32312 2632
rect 32306 2592 32312 2604
rect 32364 2592 32370 2644
rect 33134 2632 33140 2644
rect 33095 2604 33140 2632
rect 33134 2592 33140 2604
rect 33192 2592 33198 2644
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 8352 2536 10456 2564
rect 8352 2524 8358 2536
rect 4295 2468 8248 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 9272 2468 9413 2496
rect 9272 2456 9278 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 3142 2428 3148 2440
rect 3103 2400 3148 2428
rect 2041 2391 2099 2397
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 3973 2391 4031 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7248 2400 7757 2428
rect 7248 2388 7254 2400
rect 7745 2397 7757 2400
rect 7791 2428 7803 2431
rect 8202 2428 8208 2440
rect 7791 2400 8208 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 4614 2320 4620 2372
rect 4672 2360 4678 2372
rect 8404 2360 8432 2391
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 10428 2437 10456 2536
rect 15838 2524 15844 2576
rect 15896 2564 15902 2576
rect 15896 2536 18276 2564
rect 15896 2524 15902 2536
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11756 2468 11989 2496
rect 11756 2456 11762 2468
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12253 2499 12311 2505
rect 12253 2465 12265 2499
rect 12299 2496 12311 2499
rect 13538 2496 13544 2508
rect 12299 2468 13544 2496
rect 12299 2465 12311 2468
rect 12253 2459 12311 2465
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 14752 2468 15976 2496
rect 14752 2437 14780 2468
rect 15948 2440 15976 2468
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8536 2400 9137 2428
rect 8536 2388 8542 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 15378 2428 15384 2440
rect 15339 2400 15384 2428
rect 14737 2391 14795 2397
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15988 2400 16037 2428
rect 15988 2388 15994 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17000 2400 17509 2428
rect 17000 2388 17006 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2397 18199 2431
rect 18248 2428 18276 2536
rect 19426 2524 19432 2576
rect 19484 2564 19490 2576
rect 20717 2567 20775 2573
rect 20717 2564 20729 2567
rect 19484 2536 20729 2564
rect 19484 2524 19490 2536
rect 20717 2533 20729 2536
rect 20763 2533 20775 2567
rect 23474 2564 23480 2576
rect 20717 2527 20775 2533
rect 20824 2536 23480 2564
rect 19242 2456 19248 2508
rect 19300 2496 19306 2508
rect 20824 2496 20852 2536
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 19300 2468 20852 2496
rect 19300 2456 19306 2468
rect 21818 2456 21824 2508
rect 21876 2496 21882 2508
rect 21876 2468 22692 2496
rect 21876 2456 21882 2468
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 18248 2400 19441 2428
rect 18141 2391 18199 2397
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 19429 2391 19487 2397
rect 8570 2360 8576 2372
rect 4672 2332 8576 2360
rect 4672 2320 4678 2332
rect 8570 2320 8576 2332
rect 8628 2320 8634 2372
rect 9950 2320 9956 2372
rect 10008 2360 10014 2372
rect 10502 2360 10508 2372
rect 10008 2332 10508 2360
rect 10008 2320 10014 2332
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 17954 2360 17960 2372
rect 13478 2332 17960 2360
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 18156 2360 18184 2391
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20680 2400 20913 2428
rect 20680 2388 20686 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22664 2437 22692 2468
rect 31110 2456 31116 2508
rect 31168 2496 31174 2508
rect 31168 2468 35894 2496
rect 31168 2456 31174 2468
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21968 2400 22201 2428
rect 21968 2388 21974 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 23566 2428 23572 2440
rect 23527 2400 23572 2428
rect 22649 2391 22707 2397
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 23900 2400 24777 2428
rect 23900 2388 23906 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 25225 2431 25283 2437
rect 25225 2397 25237 2431
rect 25271 2428 25283 2431
rect 25590 2428 25596 2440
rect 25271 2400 25596 2428
rect 25271 2397 25283 2400
rect 25225 2391 25283 2397
rect 25590 2388 25596 2400
rect 25648 2388 25654 2440
rect 25958 2428 25964 2440
rect 25919 2400 25964 2428
rect 25958 2388 25964 2400
rect 26016 2388 26022 2440
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 29730 2428 29736 2440
rect 29691 2400 29736 2428
rect 28629 2391 28687 2397
rect 29730 2388 29736 2400
rect 29788 2388 29794 2440
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 30340 2400 30665 2428
rect 30340 2388 30346 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31570 2388 31576 2440
rect 31628 2428 31634 2440
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 31628 2400 32505 2428
rect 31628 2388 31634 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 33686 2428 33692 2440
rect 33647 2400 33692 2428
rect 32493 2391 32551 2397
rect 33686 2388 33692 2400
rect 33744 2388 33750 2440
rect 34422 2388 34428 2440
rect 34480 2428 34486 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34480 2400 34897 2428
rect 34480 2388 34486 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 35866 2428 35894 2468
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35866 2400 36185 2428
rect 34885 2391 34943 2397
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 36173 2391 36231 2397
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36780 2400 37473 2428
rect 36780 2388 36786 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37734 2428 37740 2440
rect 37695 2400 37740 2428
rect 37461 2391 37519 2397
rect 37734 2388 37740 2400
rect 37792 2388 37798 2440
rect 23290 2360 23296 2372
rect 18156 2332 23296 2360
rect 23290 2320 23296 2332
rect 23348 2320 23354 2372
rect 32858 2320 32864 2372
rect 32916 2360 32922 2372
rect 33045 2363 33103 2369
rect 33045 2360 33057 2363
rect 32916 2332 33057 2360
rect 32916 2320 32922 2332
rect 33045 2329 33057 2332
rect 33091 2329 33103 2363
rect 33045 2323 33103 2329
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 2004 2264 2237 2292
rect 2004 2252 2010 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3292 2264 3341 2292
rect 3292 2252 3298 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 8481 2295 8539 2301
rect 8481 2261 8493 2295
rect 8527 2292 8539 2295
rect 13078 2292 13084 2304
rect 8527 2264 13084 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 15470 2292 15476 2304
rect 15431 2264 15476 2292
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 19521 2295 19579 2301
rect 19521 2261 19533 2295
rect 19567 2292 19579 2295
rect 20990 2292 20996 2304
rect 19567 2264 20996 2292
rect 19567 2261 19579 2264
rect 19521 2255 19579 2261
rect 20990 2252 20996 2264
rect 21048 2252 21054 2304
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 23382 2292 23388 2304
rect 23343 2264 23388 2292
rect 22833 2255 22891 2261
rect 23382 2252 23388 2264
rect 23440 2252 23446 2304
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26145 2295 26203 2301
rect 26145 2292 26157 2295
rect 25832 2264 26157 2292
rect 25832 2252 25838 2264
rect 26145 2261 26157 2264
rect 26191 2261 26203 2295
rect 26145 2255 26203 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29696 2264 29929 2292
rect 29696 2252 29702 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33873 2295 33931 2301
rect 33873 2292 33885 2295
rect 33560 2264 33885 2292
rect 33560 2252 33566 2264
rect 33873 2261 33885 2264
rect 33919 2261 33931 2295
rect 33873 2255 33931 2261
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 36136 2264 36369 2292
rect 36136 2252 36142 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 10870 2048 10876 2100
rect 10928 2088 10934 2100
rect 27246 2088 27252 2100
rect 10928 2060 27252 2088
rect 10928 2048 10934 2060
rect 27246 2048 27252 2060
rect 27304 2048 27310 2100
rect 3602 1980 3608 2032
rect 3660 2020 3666 2032
rect 15470 2020 15476 2032
rect 3660 1992 15476 2020
rect 3660 1980 3666 1992
rect 15470 1980 15476 1992
rect 15528 1980 15534 2032
rect 17954 1980 17960 2032
rect 18012 2020 18018 2032
rect 24854 2020 24860 2032
rect 18012 1992 24860 2020
rect 18012 1980 18018 1992
rect 24854 1980 24860 1992
rect 24912 1980 24918 2032
rect 10778 1912 10784 1964
rect 10836 1952 10842 1964
rect 10836 1924 20024 1952
rect 10836 1912 10842 1924
rect 9030 1844 9036 1896
rect 9088 1884 9094 1896
rect 19242 1884 19248 1896
rect 9088 1856 19248 1884
rect 9088 1844 9094 1856
rect 19242 1844 19248 1856
rect 19300 1844 19306 1896
rect 19996 1884 20024 1924
rect 20070 1912 20076 1964
rect 20128 1952 20134 1964
rect 26694 1952 26700 1964
rect 20128 1924 26700 1952
rect 20128 1912 20134 1924
rect 26694 1912 26700 1924
rect 26752 1912 26758 1964
rect 24118 1884 24124 1896
rect 19996 1856 24124 1884
rect 24118 1844 24124 1856
rect 24176 1844 24182 1896
rect 8570 1776 8576 1828
rect 8628 1816 8634 1828
rect 15378 1816 15384 1828
rect 8628 1788 15384 1816
rect 8628 1776 8634 1788
rect 15378 1776 15384 1788
rect 15436 1776 15442 1828
rect 37734 1816 37740 1828
rect 26206 1788 37740 1816
rect 13722 1708 13728 1760
rect 13780 1748 13786 1760
rect 22186 1748 22192 1760
rect 13780 1720 22192 1748
rect 13780 1708 13786 1720
rect 22186 1708 22192 1720
rect 22244 1708 22250 1760
rect 22278 1708 22284 1760
rect 22336 1748 22342 1760
rect 26206 1748 26234 1788
rect 37734 1776 37740 1788
rect 37792 1776 37798 1828
rect 22336 1720 26234 1748
rect 22336 1708 22342 1720
rect 16114 1640 16120 1692
rect 16172 1680 16178 1692
rect 17310 1680 17316 1692
rect 16172 1652 17316 1680
rect 16172 1640 16178 1652
rect 17310 1640 17316 1652
rect 17368 1640 17374 1692
rect 17402 1640 17408 1692
rect 17460 1680 17466 1692
rect 23566 1680 23572 1692
rect 17460 1652 23572 1680
rect 17460 1640 17466 1652
rect 23566 1640 23572 1652
rect 23624 1640 23630 1692
rect 13814 1572 13820 1624
rect 13872 1612 13878 1624
rect 21542 1612 21548 1624
rect 13872 1584 21548 1612
rect 13872 1572 13878 1584
rect 21542 1572 21548 1584
rect 21600 1572 21606 1624
rect 20530 1300 20536 1352
rect 20588 1340 20594 1352
rect 25682 1340 25688 1352
rect 20588 1312 25688 1340
rect 20588 1300 20594 1312
rect 25682 1300 25688 1312
rect 25740 1300 25746 1352
rect 14826 1232 14832 1284
rect 14884 1272 14890 1284
rect 24762 1272 24768 1284
rect 14884 1244 24768 1272
rect 14884 1232 14890 1244
rect 24762 1232 24768 1244
rect 24820 1232 24826 1284
rect 4982 1164 4988 1216
rect 5040 1204 5046 1216
rect 21266 1204 21272 1216
rect 5040 1176 21272 1204
rect 5040 1164 5046 1176
rect 21266 1164 21272 1176
rect 21324 1164 21330 1216
rect 10870 144 10876 196
rect 10928 184 10934 196
rect 24946 184 24952 196
rect 10928 156 24952 184
rect 10928 144 10934 156
rect 24946 144 24952 156
rect 25004 144 25010 196
rect 11698 76 11704 128
rect 11756 116 11762 128
rect 27982 116 27988 128
rect 11756 88 27988 116
rect 11756 76 11762 88
rect 27982 76 27988 88
rect 28040 76 28046 128
rect 7190 8 7196 60
rect 7248 48 7254 60
rect 27338 48 27344 60
rect 7248 20 27344 48
rect 7248 8 7254 20
rect 27338 8 27344 20
rect 27396 8 27402 60
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1584 37315 1636 37324
rect 1584 37281 1593 37315
rect 1593 37281 1627 37315
rect 1627 37281 1636 37315
rect 1584 37272 1636 37281
rect 2872 37247 2924 37256
rect 2872 37213 2881 37247
rect 2881 37213 2915 37247
rect 2915 37213 2924 37247
rect 2872 37204 2924 37213
rect 3240 37204 3292 37256
rect 4620 37204 4672 37256
rect 10968 37272 11020 37324
rect 21272 37272 21324 37324
rect 30932 37315 30984 37324
rect 30932 37281 30941 37315
rect 30941 37281 30975 37315
rect 30975 37281 30984 37315
rect 30932 37272 30984 37281
rect 34152 37272 34204 37324
rect 38660 37272 38712 37324
rect 5540 37204 5592 37256
rect 5816 37204 5868 37256
rect 6460 37204 6512 37256
rect 7840 37247 7892 37256
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 9772 37247 9824 37256
rect 9772 37213 9781 37247
rect 9781 37213 9815 37247
rect 9815 37213 9824 37247
rect 9772 37204 9824 37213
rect 11796 37204 11848 37256
rect 12440 37204 12492 37256
rect 14280 37247 14332 37256
rect 14280 37213 14289 37247
rect 14289 37213 14323 37247
rect 14323 37213 14332 37247
rect 14280 37204 14332 37213
rect 15476 37204 15528 37256
rect 17500 37247 17552 37256
rect 17500 37213 17509 37247
rect 17509 37213 17543 37247
rect 17543 37213 17552 37247
rect 17500 37204 17552 37213
rect 19432 37204 19484 37256
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 24584 37247 24636 37256
rect 2780 37068 2832 37120
rect 3976 37111 4028 37120
rect 3976 37077 3985 37111
rect 3985 37077 4019 37111
rect 4019 37077 4028 37111
rect 3976 37068 4028 37077
rect 9404 37136 9456 37188
rect 18788 37136 18840 37188
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 25136 37204 25188 37256
rect 26424 37204 26476 37256
rect 27804 37247 27856 37256
rect 27804 37213 27813 37247
rect 27813 37213 27847 37247
rect 27847 37213 27856 37247
rect 27804 37204 27856 37213
rect 28356 37204 28408 37256
rect 29644 37204 29696 37256
rect 32312 37247 32364 37256
rect 22376 37136 22428 37188
rect 32312 37213 32321 37247
rect 32321 37213 32355 37247
rect 32355 37213 32364 37247
rect 32312 37204 32364 37213
rect 32864 37204 32916 37256
rect 35440 37204 35492 37256
rect 35992 37204 36044 37256
rect 31300 37136 31352 37188
rect 5816 37111 5868 37120
rect 5816 37077 5825 37111
rect 5825 37077 5859 37111
rect 5859 37077 5868 37111
rect 5816 37068 5868 37077
rect 6552 37111 6604 37120
rect 6552 37077 6561 37111
rect 6561 37077 6595 37111
rect 6595 37077 6604 37111
rect 6552 37068 6604 37077
rect 7748 37068 7800 37120
rect 9680 37068 9732 37120
rect 12348 37068 12400 37120
rect 13544 37068 13596 37120
rect 15568 37111 15620 37120
rect 15568 37077 15577 37111
rect 15577 37077 15611 37111
rect 15611 37077 15620 37111
rect 15568 37068 15620 37077
rect 17408 37068 17460 37120
rect 19340 37068 19392 37120
rect 19984 37068 20036 37120
rect 24492 37068 24544 37120
rect 25320 37111 25372 37120
rect 25320 37077 25329 37111
rect 25329 37077 25363 37111
rect 25363 37077 25372 37111
rect 25320 37068 25372 37077
rect 27160 37111 27212 37120
rect 27160 37077 27169 37111
rect 27169 37077 27203 37111
rect 27203 37077 27212 37111
rect 27160 37068 27212 37077
rect 27712 37068 27764 37120
rect 28540 37111 28592 37120
rect 28540 37077 28549 37111
rect 28549 37077 28583 37111
rect 28583 37077 28592 37111
rect 28540 37068 28592 37077
rect 28632 37068 28684 37120
rect 32220 37068 32272 37120
rect 33048 37111 33100 37120
rect 33048 37077 33057 37111
rect 33057 37077 33091 37111
rect 33091 37077 33100 37111
rect 33048 37068 33100 37077
rect 35532 37068 35584 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 9036 36864 9088 36916
rect 14280 36864 14332 36916
rect 16764 36864 16816 36916
rect 22100 36864 22152 36916
rect 27804 36864 27856 36916
rect 39304 36864 39356 36916
rect 1308 36796 1360 36848
rect 20 36728 72 36780
rect 14188 36796 14240 36848
rect 9128 36771 9180 36780
rect 9128 36737 9137 36771
rect 9137 36737 9171 36771
rect 9171 36737 9180 36771
rect 9128 36728 9180 36737
rect 13544 36728 13596 36780
rect 19156 36796 19208 36848
rect 22376 36796 22428 36848
rect 1860 36703 1912 36712
rect 1860 36669 1869 36703
rect 1869 36669 1903 36703
rect 1903 36669 1912 36703
rect 1860 36660 1912 36669
rect 15384 36728 15436 36780
rect 18052 36728 18104 36780
rect 23204 36728 23256 36780
rect 26240 36771 26292 36780
rect 26240 36737 26249 36771
rect 26249 36737 26283 36771
rect 26283 36737 26292 36771
rect 26240 36728 26292 36737
rect 31300 36728 31352 36780
rect 36084 36796 36136 36848
rect 38108 36839 38160 36848
rect 38108 36805 38117 36839
rect 38117 36805 38151 36839
rect 38151 36805 38160 36839
rect 38108 36796 38160 36805
rect 36176 36771 36228 36780
rect 36176 36737 36185 36771
rect 36185 36737 36219 36771
rect 36219 36737 36228 36771
rect 36176 36728 36228 36737
rect 20628 36660 20680 36712
rect 5724 36524 5776 36576
rect 33140 36524 33192 36576
rect 37924 36524 37976 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1768 36363 1820 36372
rect 1768 36329 1777 36363
rect 1777 36329 1811 36363
rect 1811 36329 1820 36363
rect 1768 36320 1820 36329
rect 9128 36320 9180 36372
rect 18604 36320 18656 36372
rect 36176 36320 36228 36372
rect 37188 36320 37240 36372
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 2780 36116 2832 36168
rect 35532 36159 35584 36168
rect 35532 36125 35541 36159
rect 35541 36125 35575 36159
rect 35575 36125 35584 36159
rect 35532 36116 35584 36125
rect 36820 36159 36872 36168
rect 36820 36125 36829 36159
rect 36829 36125 36863 36159
rect 36863 36125 36872 36159
rect 36820 36116 36872 36125
rect 37280 36159 37332 36168
rect 37280 36125 37289 36159
rect 37289 36125 37323 36159
rect 37323 36125 37332 36159
rect 37280 36116 37332 36125
rect 6828 35980 6880 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 18696 35776 18748 35828
rect 19432 35776 19484 35828
rect 4620 35640 4672 35692
rect 37832 35640 37884 35692
rect 1768 35479 1820 35488
rect 1768 35445 1777 35479
rect 1777 35445 1811 35479
rect 1811 35445 1820 35479
rect 1768 35436 1820 35445
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 22284 35164 22336 35216
rect 37280 35164 37332 35216
rect 1768 35071 1820 35080
rect 1768 35037 1777 35071
rect 1777 35037 1811 35071
rect 1811 35037 1820 35071
rect 1768 35028 1820 35037
rect 37372 35028 37424 35080
rect 4068 34892 4120 34944
rect 37464 34935 37516 34944
rect 37464 34901 37473 34935
rect 37473 34901 37507 34935
rect 37507 34901 37516 34935
rect 37464 34892 37516 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 15384 34688 15436 34740
rect 36820 34688 36872 34740
rect 13912 34552 13964 34604
rect 35440 34595 35492 34604
rect 35440 34561 35449 34595
rect 35449 34561 35483 34595
rect 35483 34561 35492 34595
rect 35440 34552 35492 34561
rect 35992 34552 36044 34604
rect 21364 34484 21416 34536
rect 24584 34484 24636 34536
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 19156 33507 19208 33516
rect 19156 33473 19165 33507
rect 19165 33473 19199 33507
rect 19199 33473 19208 33507
rect 19156 33464 19208 33473
rect 1768 33371 1820 33380
rect 1768 33337 1777 33371
rect 1777 33337 1811 33371
rect 1811 33337 1820 33371
rect 1768 33328 1820 33337
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 5724 32895 5776 32904
rect 5724 32861 5733 32895
rect 5733 32861 5767 32895
rect 5767 32861 5776 32895
rect 5724 32852 5776 32861
rect 28540 32852 28592 32904
rect 36452 32852 36504 32904
rect 6644 32716 6696 32768
rect 17776 32716 17828 32768
rect 38200 32759 38252 32768
rect 38200 32725 38209 32759
rect 38209 32725 38243 32759
rect 38243 32725 38252 32759
rect 38200 32716 38252 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 5816 32376 5868 32428
rect 33232 32376 33284 32428
rect 1584 32351 1636 32360
rect 1584 32317 1593 32351
rect 1593 32317 1627 32351
rect 1627 32317 1636 32351
rect 1584 32308 1636 32317
rect 9312 32308 9364 32360
rect 9128 32215 9180 32224
rect 9128 32181 9137 32215
rect 9137 32181 9171 32215
rect 9171 32181 9180 32215
rect 9128 32172 9180 32181
rect 38200 32215 38252 32224
rect 38200 32181 38209 32215
rect 38209 32181 38243 32215
rect 38243 32181 38252 32215
rect 38200 32172 38252 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4620 31968 4672 32020
rect 7840 31968 7892 32020
rect 17408 31968 17460 32020
rect 9036 31900 9088 31952
rect 20260 31900 20312 31952
rect 6552 31832 6604 31884
rect 4620 31764 4672 31816
rect 6736 31764 6788 31816
rect 7656 31807 7708 31816
rect 7656 31773 7665 31807
rect 7665 31773 7699 31807
rect 7699 31773 7708 31807
rect 7656 31764 7708 31773
rect 14188 31832 14240 31884
rect 19340 31764 19392 31816
rect 25320 31832 25372 31884
rect 28632 31764 28684 31816
rect 1768 31671 1820 31680
rect 1768 31637 1777 31671
rect 1777 31637 1811 31671
rect 1811 31637 1820 31671
rect 1768 31628 1820 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 7656 31424 7708 31476
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 26240 31288 26292 31340
rect 37464 31288 37516 31340
rect 20352 31084 20404 31136
rect 26700 31084 26752 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4068 30676 4120 30728
rect 9404 30719 9456 30728
rect 9404 30685 9413 30719
rect 9413 30685 9447 30719
rect 9447 30685 9456 30719
rect 9404 30676 9456 30685
rect 27160 30676 27212 30728
rect 38292 30719 38344 30728
rect 38292 30685 38301 30719
rect 38301 30685 38335 30719
rect 38335 30685 38344 30719
rect 38292 30676 38344 30685
rect 1860 30608 1912 30660
rect 33692 30608 33744 30660
rect 8576 30540 8628 30592
rect 11336 30540 11388 30592
rect 17132 30540 17184 30592
rect 37004 30540 37056 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 5448 30200 5500 30252
rect 12348 30243 12400 30252
rect 12348 30209 12357 30243
rect 12357 30209 12391 30243
rect 12391 30209 12400 30243
rect 12348 30200 12400 30209
rect 33048 30268 33100 30320
rect 33140 30200 33192 30252
rect 17224 30064 17276 30116
rect 1768 30039 1820 30048
rect 1768 30005 1777 30039
rect 1777 30005 1811 30039
rect 1811 30005 1820 30039
rect 1768 29996 1820 30005
rect 12440 30039 12492 30048
rect 12440 30005 12449 30039
rect 12449 30005 12483 30039
rect 12483 30005 12492 30039
rect 12440 29996 12492 30005
rect 18236 29996 18288 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 6736 29835 6788 29844
rect 6736 29801 6745 29835
rect 6745 29801 6779 29835
rect 6779 29801 6788 29835
rect 6736 29792 6788 29801
rect 3976 29656 4028 29708
rect 8944 29588 8996 29640
rect 19984 29588 20036 29640
rect 35900 29588 35952 29640
rect 38108 29563 38160 29572
rect 38108 29529 38117 29563
rect 38117 29529 38151 29563
rect 38151 29529 38160 29563
rect 38108 29520 38160 29529
rect 10600 29452 10652 29504
rect 37740 29452 37792 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4620 29248 4672 29300
rect 33232 29291 33284 29300
rect 33232 29257 33241 29291
rect 33241 29257 33275 29291
rect 33275 29257 33284 29291
rect 33232 29248 33284 29257
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 5908 29112 5960 29164
rect 6828 29112 6880 29164
rect 31760 29112 31812 29164
rect 2688 28976 2740 29028
rect 6828 28976 6880 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 15568 28500 15620 28552
rect 35440 28500 35492 28552
rect 2872 28432 2924 28484
rect 20720 28432 20772 28484
rect 15752 28364 15804 28416
rect 24860 28364 24912 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 36452 28160 36504 28212
rect 15200 28092 15252 28144
rect 1400 28024 1452 28076
rect 19156 28024 19208 28076
rect 24032 28024 24084 28076
rect 38292 28067 38344 28076
rect 38292 28033 38301 28067
rect 38301 28033 38335 28067
rect 38335 28033 38344 28067
rect 38292 28024 38344 28033
rect 17960 27888 18012 27940
rect 5172 27820 5224 27872
rect 11244 27820 11296 27872
rect 14188 27820 14240 27872
rect 18144 27820 18196 27872
rect 36084 27820 36136 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 31760 27548 31812 27600
rect 6000 27480 6052 27532
rect 12348 27480 12400 27532
rect 2412 27412 2464 27464
rect 11980 27412 12032 27464
rect 13544 27455 13596 27464
rect 13544 27421 13553 27455
rect 13553 27421 13587 27455
rect 13587 27421 13596 27455
rect 13544 27412 13596 27421
rect 13636 27412 13688 27464
rect 26240 27412 26292 27464
rect 35900 27412 35952 27464
rect 5264 27344 5316 27396
rect 9772 27344 9824 27396
rect 14464 27344 14516 27396
rect 1768 27319 1820 27328
rect 1768 27285 1777 27319
rect 1777 27285 1811 27319
rect 1811 27285 1820 27319
rect 1768 27276 1820 27285
rect 2504 27276 2556 27328
rect 11060 27276 11112 27328
rect 12256 27319 12308 27328
rect 12256 27285 12265 27319
rect 12265 27285 12299 27319
rect 12299 27285 12308 27319
rect 12256 27276 12308 27285
rect 12624 27276 12676 27328
rect 13452 27276 13504 27328
rect 14372 27319 14424 27328
rect 14372 27285 14381 27319
rect 14381 27285 14415 27319
rect 14415 27285 14424 27319
rect 14372 27276 14424 27285
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 5908 27115 5960 27124
rect 5908 27081 5917 27115
rect 5917 27081 5951 27115
rect 5951 27081 5960 27115
rect 5908 27072 5960 27081
rect 8208 27072 8260 27124
rect 8944 27004 8996 27056
rect 1860 26979 1912 26988
rect 1860 26945 1869 26979
rect 1869 26945 1903 26979
rect 1903 26945 1912 26979
rect 1860 26936 1912 26945
rect 2320 26936 2372 26988
rect 5816 26979 5868 26988
rect 5816 26945 5825 26979
rect 5825 26945 5859 26979
rect 5859 26945 5868 26979
rect 5816 26936 5868 26945
rect 6460 26936 6512 26988
rect 11060 26979 11112 26988
rect 7840 26868 7892 26920
rect 6736 26800 6788 26852
rect 11060 26945 11069 26979
rect 11069 26945 11103 26979
rect 11103 26945 11112 26979
rect 11060 26936 11112 26945
rect 15200 27072 15252 27124
rect 14372 27004 14424 27056
rect 12348 26979 12400 26988
rect 12348 26945 12357 26979
rect 12357 26945 12391 26979
rect 12391 26945 12400 26979
rect 12348 26936 12400 26945
rect 14464 26979 14516 26988
rect 14464 26945 14473 26979
rect 14473 26945 14507 26979
rect 14507 26945 14516 26979
rect 14464 26936 14516 26945
rect 37004 26936 37056 26988
rect 10876 26868 10928 26920
rect 10968 26868 11020 26920
rect 14004 26868 14056 26920
rect 1676 26732 1728 26784
rect 2596 26775 2648 26784
rect 2596 26741 2605 26775
rect 2605 26741 2639 26775
rect 2639 26741 2648 26775
rect 2596 26732 2648 26741
rect 3240 26775 3292 26784
rect 3240 26741 3249 26775
rect 3249 26741 3283 26775
rect 3283 26741 3292 26775
rect 3240 26732 3292 26741
rect 8024 26775 8076 26784
rect 8024 26741 8033 26775
rect 8033 26741 8067 26775
rect 8067 26741 8076 26775
rect 8024 26732 8076 26741
rect 10048 26732 10100 26784
rect 13820 26800 13872 26852
rect 13912 26843 13964 26852
rect 13912 26809 13921 26843
rect 13921 26809 13955 26843
rect 13955 26809 13964 26843
rect 13912 26800 13964 26809
rect 11980 26732 12032 26784
rect 12532 26732 12584 26784
rect 32404 26775 32456 26784
rect 32404 26741 32413 26775
rect 32413 26741 32447 26775
rect 32447 26741 32456 26775
rect 32404 26732 32456 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 18052 26571 18104 26580
rect 4068 26460 4120 26512
rect 9312 26460 9364 26512
rect 10140 26460 10192 26512
rect 10876 26460 10928 26512
rect 11888 26460 11940 26512
rect 2228 26324 2280 26376
rect 2688 26367 2740 26376
rect 2688 26333 2697 26367
rect 2697 26333 2731 26367
rect 2731 26333 2740 26367
rect 2688 26324 2740 26333
rect 4804 26324 4856 26376
rect 6460 26367 6512 26376
rect 6460 26333 6469 26367
rect 6469 26333 6503 26367
rect 6503 26333 6512 26367
rect 6460 26324 6512 26333
rect 10048 26435 10100 26444
rect 10048 26401 10057 26435
rect 10057 26401 10091 26435
rect 10091 26401 10100 26435
rect 10048 26392 10100 26401
rect 10968 26435 11020 26444
rect 10968 26401 10977 26435
rect 10977 26401 11011 26435
rect 11011 26401 11020 26435
rect 10968 26392 11020 26401
rect 13912 26392 13964 26444
rect 11152 26367 11204 26376
rect 11152 26333 11161 26367
rect 11161 26333 11195 26367
rect 11195 26333 11204 26367
rect 11152 26324 11204 26333
rect 12256 26367 12308 26376
rect 12256 26333 12265 26367
rect 12265 26333 12299 26367
rect 12299 26333 12308 26367
rect 12256 26324 12308 26333
rect 18052 26537 18061 26571
rect 18061 26537 18095 26571
rect 18095 26537 18104 26571
rect 18052 26528 18104 26537
rect 19064 26460 19116 26512
rect 35992 26528 36044 26580
rect 34612 26460 34664 26512
rect 24860 26392 24912 26444
rect 17592 26324 17644 26376
rect 19340 26324 19392 26376
rect 38292 26367 38344 26376
rect 2320 26256 2372 26308
rect 2964 26256 3016 26308
rect 9588 26256 9640 26308
rect 11152 26188 11204 26240
rect 16396 26256 16448 26308
rect 17316 26256 17368 26308
rect 20168 26256 20220 26308
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 19432 26231 19484 26240
rect 19432 26197 19441 26231
rect 19441 26197 19475 26231
rect 19475 26197 19484 26231
rect 19432 26188 19484 26197
rect 22836 26231 22888 26240
rect 22836 26197 22845 26231
rect 22845 26197 22879 26231
rect 22879 26197 22888 26231
rect 22836 26188 22888 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 9220 25984 9272 26036
rect 1124 25848 1176 25900
rect 1216 25780 1268 25832
rect 4896 25891 4948 25900
rect 2872 25780 2924 25832
rect 4896 25857 4905 25891
rect 4905 25857 4939 25891
rect 4939 25857 4948 25891
rect 4896 25848 4948 25857
rect 7012 25780 7064 25832
rect 7196 25780 7248 25832
rect 14004 25984 14056 26036
rect 18604 25984 18656 26036
rect 20444 25984 20496 26036
rect 8024 25891 8076 25900
rect 8024 25857 8033 25891
rect 8033 25857 8067 25891
rect 8067 25857 8076 25891
rect 8024 25848 8076 25857
rect 9404 25891 9456 25900
rect 9404 25857 9413 25891
rect 9413 25857 9447 25891
rect 9447 25857 9456 25891
rect 9404 25848 9456 25857
rect 10784 25891 10836 25900
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 12900 25848 12952 25900
rect 18788 25916 18840 25968
rect 7932 25780 7984 25832
rect 19432 25848 19484 25900
rect 19248 25780 19300 25832
rect 6736 25712 6788 25764
rect 15936 25712 15988 25764
rect 18972 25712 19024 25764
rect 1860 25644 1912 25696
rect 3792 25644 3844 25696
rect 3976 25644 4028 25696
rect 4712 25687 4764 25696
rect 4712 25653 4721 25687
rect 4721 25653 4755 25687
rect 4755 25653 4764 25687
rect 4712 25644 4764 25653
rect 8300 25687 8352 25696
rect 8300 25653 8309 25687
rect 8309 25653 8343 25687
rect 8343 25653 8352 25687
rect 8300 25644 8352 25653
rect 10140 25644 10192 25696
rect 10232 25644 10284 25696
rect 11428 25644 11480 25696
rect 14096 25644 14148 25696
rect 18788 25687 18840 25696
rect 18788 25653 18797 25687
rect 18797 25653 18831 25687
rect 18831 25653 18840 25687
rect 18788 25644 18840 25653
rect 19340 25687 19392 25696
rect 19340 25653 19349 25687
rect 19349 25653 19383 25687
rect 19383 25653 19392 25687
rect 19340 25644 19392 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5264 25483 5316 25492
rect 5264 25449 5273 25483
rect 5273 25449 5307 25483
rect 5307 25449 5316 25483
rect 5264 25440 5316 25449
rect 11888 25440 11940 25492
rect 12900 25440 12952 25492
rect 17868 25440 17920 25492
rect 18788 25440 18840 25492
rect 31116 25440 31168 25492
rect 35900 25440 35952 25492
rect 10784 25372 10836 25424
rect 7932 25304 7984 25356
rect 11336 25347 11388 25356
rect 11336 25313 11345 25347
rect 11345 25313 11379 25347
rect 11379 25313 11388 25347
rect 11336 25304 11388 25313
rect 12532 25304 12584 25356
rect 12808 25304 12860 25356
rect 14924 25304 14976 25356
rect 17132 25347 17184 25356
rect 17132 25313 17141 25347
rect 17141 25313 17175 25347
rect 17175 25313 17184 25347
rect 17132 25304 17184 25313
rect 17500 25347 17552 25356
rect 17500 25313 17509 25347
rect 17509 25313 17543 25347
rect 17543 25313 17552 25347
rect 17500 25304 17552 25313
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 1032 25168 1084 25220
rect 3976 25279 4028 25288
rect 3976 25245 3985 25279
rect 3985 25245 4019 25279
rect 4019 25245 4028 25279
rect 3976 25236 4028 25245
rect 4528 25236 4580 25288
rect 5356 25236 5408 25288
rect 8484 25236 8536 25288
rect 9220 25236 9272 25288
rect 10784 25168 10836 25220
rect 3240 25100 3292 25152
rect 4620 25100 4672 25152
rect 6736 25100 6788 25152
rect 9680 25143 9732 25152
rect 9680 25109 9689 25143
rect 9689 25109 9723 25143
rect 9723 25109 9732 25143
rect 9680 25100 9732 25109
rect 10140 25100 10192 25152
rect 13728 25236 13780 25288
rect 19984 25372 20036 25424
rect 22836 25304 22888 25356
rect 18420 25236 18472 25288
rect 19248 25236 19300 25288
rect 24124 25236 24176 25288
rect 11428 25211 11480 25220
rect 11428 25177 11437 25211
rect 11437 25177 11471 25211
rect 11471 25177 11480 25211
rect 11428 25168 11480 25177
rect 12072 25168 12124 25220
rect 12900 25100 12952 25152
rect 16948 25100 17000 25152
rect 21916 25100 21968 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1952 24828 2004 24880
rect 2504 24828 2556 24880
rect 2688 24803 2740 24812
rect 2688 24769 2697 24803
rect 2697 24769 2731 24803
rect 2731 24769 2740 24803
rect 2688 24760 2740 24769
rect 3424 24760 3476 24812
rect 3700 24760 3752 24812
rect 4528 24760 4580 24812
rect 5632 24828 5684 24880
rect 6736 24871 6788 24880
rect 6736 24837 6745 24871
rect 6745 24837 6779 24871
rect 6779 24837 6788 24871
rect 6736 24828 6788 24837
rect 12072 24896 12124 24948
rect 17500 24896 17552 24948
rect 8116 24871 8168 24880
rect 8116 24837 8125 24871
rect 8125 24837 8159 24871
rect 8159 24837 8168 24871
rect 8116 24828 8168 24837
rect 9312 24871 9364 24880
rect 9312 24837 9321 24871
rect 9321 24837 9355 24871
rect 9355 24837 9364 24871
rect 9312 24828 9364 24837
rect 14096 24871 14148 24880
rect 5540 24760 5592 24812
rect 6552 24760 6604 24812
rect 10968 24760 11020 24812
rect 6184 24692 6236 24744
rect 8208 24692 8260 24744
rect 9220 24735 9272 24744
rect 9220 24701 9229 24735
rect 9229 24701 9263 24735
rect 9263 24701 9272 24735
rect 9220 24692 9272 24701
rect 9404 24692 9456 24744
rect 14096 24837 14105 24871
rect 14105 24837 14139 24871
rect 14139 24837 14148 24871
rect 14096 24828 14148 24837
rect 13820 24760 13872 24812
rect 15108 24803 15160 24812
rect 2044 24599 2096 24608
rect 2044 24565 2053 24599
rect 2053 24565 2087 24599
rect 2087 24565 2096 24599
rect 2044 24556 2096 24565
rect 2780 24599 2832 24608
rect 2780 24565 2789 24599
rect 2789 24565 2823 24599
rect 2823 24565 2832 24599
rect 2780 24556 2832 24565
rect 3056 24556 3108 24608
rect 3884 24599 3936 24608
rect 3884 24565 3893 24599
rect 3893 24565 3927 24599
rect 3927 24565 3936 24599
rect 3884 24556 3936 24565
rect 4988 24556 5040 24608
rect 5264 24556 5316 24608
rect 7932 24624 7984 24676
rect 7564 24556 7616 24608
rect 8944 24624 8996 24676
rect 11704 24624 11756 24676
rect 13176 24624 13228 24676
rect 14372 24692 14424 24744
rect 15108 24769 15117 24803
rect 15117 24769 15151 24803
rect 15151 24769 15160 24803
rect 15108 24760 15160 24769
rect 22192 24871 22244 24880
rect 22192 24837 22201 24871
rect 22201 24837 22235 24871
rect 22235 24837 22244 24871
rect 22192 24828 22244 24837
rect 18144 24760 18196 24812
rect 19340 24760 19392 24812
rect 20168 24803 20220 24812
rect 20168 24769 20177 24803
rect 20177 24769 20211 24803
rect 20211 24769 20220 24803
rect 20168 24760 20220 24769
rect 22836 24760 22888 24812
rect 16948 24735 17000 24744
rect 16948 24701 16957 24735
rect 16957 24701 16991 24735
rect 16991 24701 17000 24735
rect 16948 24692 17000 24701
rect 19432 24692 19484 24744
rect 21916 24692 21968 24744
rect 34520 24760 34572 24812
rect 35992 24692 36044 24744
rect 11888 24599 11940 24608
rect 11888 24565 11897 24599
rect 11897 24565 11931 24599
rect 11931 24565 11940 24599
rect 11888 24556 11940 24565
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 13544 24556 13596 24608
rect 14648 24624 14700 24676
rect 15200 24599 15252 24608
rect 15200 24565 15209 24599
rect 15209 24565 15243 24599
rect 15243 24565 15252 24599
rect 15200 24556 15252 24565
rect 16212 24624 16264 24676
rect 20168 24624 20220 24676
rect 20904 24624 20956 24676
rect 26240 24624 26292 24676
rect 17040 24556 17092 24608
rect 18696 24599 18748 24608
rect 18696 24565 18705 24599
rect 18705 24565 18739 24599
rect 18739 24565 18748 24599
rect 18696 24556 18748 24565
rect 22192 24556 22244 24608
rect 29092 24599 29144 24608
rect 29092 24565 29101 24599
rect 29101 24565 29135 24599
rect 29135 24565 29144 24599
rect 29092 24556 29144 24565
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 940 24352 992 24404
rect 3700 24352 3752 24404
rect 6184 24395 6236 24404
rect 6184 24361 6193 24395
rect 6193 24361 6227 24395
rect 6227 24361 6236 24395
rect 6184 24352 6236 24361
rect 7840 24352 7892 24404
rect 10508 24352 10560 24404
rect 11888 24352 11940 24404
rect 13084 24352 13136 24404
rect 13176 24352 13228 24404
rect 16212 24352 16264 24404
rect 17776 24352 17828 24404
rect 20076 24352 20128 24404
rect 3884 24284 3936 24336
rect 12716 24284 12768 24336
rect 4344 24216 4396 24268
rect 1492 24148 1544 24200
rect 2504 24191 2556 24200
rect 2504 24157 2513 24191
rect 2513 24157 2547 24191
rect 2547 24157 2556 24191
rect 2504 24148 2556 24157
rect 4712 24148 4764 24200
rect 4988 24191 5040 24200
rect 4988 24157 4997 24191
rect 4997 24157 5031 24191
rect 5031 24157 5040 24191
rect 4988 24148 5040 24157
rect 5632 24148 5684 24200
rect 6092 24191 6144 24200
rect 6092 24157 6101 24191
rect 6101 24157 6135 24191
rect 6135 24157 6144 24191
rect 6092 24148 6144 24157
rect 9220 24216 9272 24268
rect 12532 24259 12584 24268
rect 12532 24225 12541 24259
rect 12541 24225 12575 24259
rect 12575 24225 12584 24259
rect 13268 24284 13320 24336
rect 13176 24259 13228 24268
rect 12532 24216 12584 24225
rect 13176 24225 13185 24259
rect 13185 24225 13219 24259
rect 13219 24225 13228 24259
rect 13176 24216 13228 24225
rect 13544 24216 13596 24268
rect 3608 24080 3660 24132
rect 2504 24012 2556 24064
rect 3148 24055 3200 24064
rect 3148 24021 3157 24055
rect 3157 24021 3191 24055
rect 3191 24021 3200 24055
rect 3148 24012 3200 24021
rect 3332 24012 3384 24064
rect 4712 24012 4764 24064
rect 4988 24012 5040 24064
rect 7104 24055 7156 24064
rect 7104 24021 7113 24055
rect 7113 24021 7147 24055
rect 7147 24021 7156 24055
rect 7104 24012 7156 24021
rect 8300 24148 8352 24200
rect 10968 24148 11020 24200
rect 18052 24284 18104 24336
rect 20904 24327 20956 24336
rect 13820 24216 13872 24268
rect 17776 24216 17828 24268
rect 17868 24216 17920 24268
rect 9128 24080 9180 24132
rect 10232 24080 10284 24132
rect 10692 24123 10744 24132
rect 10692 24089 10701 24123
rect 10701 24089 10735 24123
rect 10735 24089 10744 24123
rect 10692 24080 10744 24089
rect 12624 24123 12676 24132
rect 12624 24089 12633 24123
rect 12633 24089 12667 24123
rect 12667 24089 12676 24123
rect 12624 24080 12676 24089
rect 12992 24080 13044 24132
rect 15108 24148 15160 24200
rect 18696 24216 18748 24268
rect 20904 24293 20913 24327
rect 20913 24293 20947 24327
rect 20947 24293 20956 24327
rect 20904 24284 20956 24293
rect 18328 24148 18380 24200
rect 19524 24148 19576 24200
rect 22836 24191 22888 24200
rect 22836 24157 22845 24191
rect 22845 24157 22879 24191
rect 22879 24157 22888 24191
rect 22836 24148 22888 24157
rect 24308 24148 24360 24200
rect 36084 24148 36136 24200
rect 9772 24012 9824 24064
rect 11244 24055 11296 24064
rect 11244 24021 11253 24055
rect 11253 24021 11287 24055
rect 11287 24021 11296 24055
rect 11244 24012 11296 24021
rect 12440 24012 12492 24064
rect 19340 24080 19392 24132
rect 14372 24055 14424 24064
rect 14372 24021 14381 24055
rect 14381 24021 14415 24055
rect 14415 24021 14424 24055
rect 14372 24012 14424 24021
rect 15016 24055 15068 24064
rect 15016 24021 15025 24055
rect 15025 24021 15059 24055
rect 15059 24021 15068 24055
rect 15016 24012 15068 24021
rect 17592 24012 17644 24064
rect 19248 24012 19300 24064
rect 38200 24055 38252 24064
rect 38200 24021 38209 24055
rect 38209 24021 38243 24055
rect 38243 24021 38252 24055
rect 38200 24012 38252 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3608 23808 3660 23860
rect 4620 23740 4672 23792
rect 1400 23672 1452 23724
rect 5172 23740 5224 23792
rect 2136 23647 2188 23656
rect 2136 23613 2145 23647
rect 2145 23613 2179 23647
rect 2179 23613 2188 23647
rect 2136 23604 2188 23613
rect 1308 23536 1360 23588
rect 3056 23536 3108 23588
rect 2044 23468 2096 23520
rect 2688 23468 2740 23520
rect 3608 23604 3660 23656
rect 5080 23672 5132 23724
rect 5448 23808 5500 23860
rect 8576 23783 8628 23792
rect 8576 23749 8585 23783
rect 8585 23749 8619 23783
rect 8619 23749 8628 23783
rect 8576 23740 8628 23749
rect 9680 23808 9732 23860
rect 5632 23715 5684 23724
rect 5632 23681 5641 23715
rect 5641 23681 5675 23715
rect 5675 23681 5684 23715
rect 5632 23672 5684 23681
rect 6460 23672 6512 23724
rect 7012 23672 7064 23724
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 9772 23672 9824 23724
rect 10324 23672 10376 23724
rect 11060 23672 11112 23724
rect 12440 23808 12492 23860
rect 15016 23808 15068 23860
rect 15108 23808 15160 23860
rect 18052 23808 18104 23860
rect 18696 23808 18748 23860
rect 19800 23808 19852 23860
rect 29092 23808 29144 23860
rect 13728 23783 13780 23792
rect 13728 23749 13737 23783
rect 13737 23749 13771 23783
rect 13771 23749 13780 23783
rect 13728 23740 13780 23749
rect 17592 23783 17644 23792
rect 17592 23749 17601 23783
rect 17601 23749 17635 23783
rect 17635 23749 17644 23783
rect 17592 23740 17644 23749
rect 17776 23740 17828 23792
rect 37740 23740 37792 23792
rect 14832 23715 14884 23724
rect 3976 23536 4028 23588
rect 5816 23604 5868 23656
rect 6184 23604 6236 23656
rect 14832 23681 14841 23715
rect 14841 23681 14875 23715
rect 14875 23681 14884 23715
rect 14832 23672 14884 23681
rect 15936 23715 15988 23724
rect 15936 23681 15945 23715
rect 15945 23681 15979 23715
rect 15979 23681 15988 23715
rect 15936 23672 15988 23681
rect 19248 23715 19300 23724
rect 19248 23681 19257 23715
rect 19257 23681 19291 23715
rect 19291 23681 19300 23715
rect 19248 23672 19300 23681
rect 20168 23672 20220 23724
rect 23480 23715 23532 23724
rect 6000 23536 6052 23588
rect 7840 23536 7892 23588
rect 12992 23604 13044 23656
rect 8668 23536 8720 23588
rect 13728 23604 13780 23656
rect 17960 23647 18012 23656
rect 13912 23536 13964 23588
rect 15660 23536 15712 23588
rect 17960 23613 17969 23647
rect 17969 23613 18003 23647
rect 18003 23613 18012 23647
rect 17960 23604 18012 23613
rect 18788 23604 18840 23656
rect 19524 23604 19576 23656
rect 20352 23604 20404 23656
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 23480 23672 23532 23681
rect 34612 23672 34664 23724
rect 24584 23604 24636 23656
rect 18236 23536 18288 23588
rect 4344 23468 4396 23520
rect 4620 23468 4672 23520
rect 5172 23468 5224 23520
rect 5632 23468 5684 23520
rect 9772 23511 9824 23520
rect 9772 23477 9781 23511
rect 9781 23477 9815 23511
rect 9815 23477 9824 23511
rect 9772 23468 9824 23477
rect 10876 23468 10928 23520
rect 12624 23468 12676 23520
rect 13084 23468 13136 23520
rect 15476 23468 15528 23520
rect 17040 23468 17092 23520
rect 19800 23468 19852 23520
rect 19984 23468 20036 23520
rect 23296 23511 23348 23520
rect 23296 23477 23305 23511
rect 23305 23477 23339 23511
rect 23339 23477 23348 23511
rect 23296 23468 23348 23477
rect 29000 23468 29052 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 6552 23264 6604 23316
rect 7932 23264 7984 23316
rect 3516 23196 3568 23248
rect 4804 23196 4856 23248
rect 2964 23128 3016 23180
rect 8852 23196 8904 23248
rect 3056 23060 3108 23112
rect 4068 23103 4120 23112
rect 4068 23069 4077 23103
rect 4077 23069 4111 23103
rect 4111 23069 4120 23103
rect 4068 23060 4120 23069
rect 5724 23060 5776 23112
rect 6368 23060 6420 23112
rect 1768 23035 1820 23044
rect 1768 23001 1777 23035
rect 1777 23001 1811 23035
rect 1811 23001 1820 23035
rect 1768 22992 1820 23001
rect 3792 22992 3844 23044
rect 6828 23060 6880 23112
rect 9496 23128 9548 23180
rect 11152 23171 11204 23180
rect 8576 23060 8628 23112
rect 6920 22992 6972 23044
rect 2596 22924 2648 22976
rect 3516 22924 3568 22976
rect 5448 22924 5500 22976
rect 5816 22924 5868 22976
rect 9680 22992 9732 23044
rect 7472 22924 7524 22976
rect 8208 22924 8260 22976
rect 9312 22967 9364 22976
rect 9312 22933 9321 22967
rect 9321 22933 9355 22967
rect 9355 22933 9364 22967
rect 9312 22924 9364 22933
rect 10048 23035 10100 23044
rect 10048 23001 10057 23035
rect 10057 23001 10091 23035
rect 10091 23001 10100 23035
rect 11152 23137 11161 23171
rect 11161 23137 11195 23171
rect 11195 23137 11204 23171
rect 11152 23128 11204 23137
rect 14740 23264 14792 23316
rect 15108 23264 15160 23316
rect 17684 23264 17736 23316
rect 34520 23264 34572 23316
rect 14372 23196 14424 23248
rect 14832 23196 14884 23248
rect 10048 22992 10100 23001
rect 13268 23128 13320 23180
rect 12532 23103 12584 23112
rect 12532 23069 12541 23103
rect 12541 23069 12575 23103
rect 12575 23069 12584 23103
rect 12532 23060 12584 23069
rect 13820 23128 13872 23180
rect 15200 23128 15252 23180
rect 17408 23128 17460 23180
rect 19524 23171 19576 23180
rect 19524 23137 19533 23171
rect 19533 23137 19567 23171
rect 19567 23137 19576 23171
rect 19524 23128 19576 23137
rect 18512 23103 18564 23112
rect 18512 23069 18521 23103
rect 18521 23069 18555 23103
rect 18555 23069 18564 23103
rect 18512 23060 18564 23069
rect 23296 23103 23348 23112
rect 23296 23069 23305 23103
rect 23305 23069 23339 23103
rect 23339 23069 23348 23103
rect 23296 23060 23348 23069
rect 12440 22924 12492 22976
rect 14096 22924 14148 22976
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 15568 22992 15620 23044
rect 15660 22924 15712 22976
rect 17132 22992 17184 23044
rect 17316 23035 17368 23044
rect 17316 23001 17325 23035
rect 17325 23001 17359 23035
rect 17359 23001 17368 23035
rect 17316 22992 17368 23001
rect 20168 23035 20220 23044
rect 16764 22924 16816 22976
rect 19340 22924 19392 22976
rect 20168 23001 20177 23035
rect 20177 23001 20211 23035
rect 20211 23001 20220 23035
rect 20168 22992 20220 23001
rect 22192 22924 22244 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 3240 22720 3292 22772
rect 8116 22720 8168 22772
rect 2780 22652 2832 22704
rect 3516 22652 3568 22704
rect 9956 22720 10008 22772
rect 10048 22720 10100 22772
rect 10140 22695 10192 22704
rect 2136 22559 2188 22568
rect 2136 22525 2145 22559
rect 2145 22525 2179 22559
rect 2179 22525 2188 22559
rect 2136 22516 2188 22525
rect 5540 22584 5592 22636
rect 5724 22584 5776 22636
rect 6000 22584 6052 22636
rect 6276 22584 6328 22636
rect 6828 22627 6880 22636
rect 6828 22593 6837 22627
rect 6837 22593 6871 22627
rect 6871 22593 6880 22627
rect 6828 22584 6880 22593
rect 8576 22584 8628 22636
rect 9128 22584 9180 22636
rect 6092 22516 6144 22568
rect 3792 22448 3844 22500
rect 10140 22661 10149 22695
rect 10149 22661 10183 22695
rect 10183 22661 10192 22695
rect 10140 22652 10192 22661
rect 10232 22652 10284 22704
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 12624 22695 12676 22704
rect 12624 22661 12633 22695
rect 12633 22661 12667 22695
rect 12667 22661 12676 22695
rect 12624 22652 12676 22661
rect 13176 22695 13228 22704
rect 13176 22661 13185 22695
rect 13185 22661 13219 22695
rect 13219 22661 13228 22695
rect 13176 22652 13228 22661
rect 14280 22720 14332 22772
rect 15476 22720 15528 22772
rect 29736 22720 29788 22772
rect 13820 22695 13872 22704
rect 13820 22661 13829 22695
rect 13829 22661 13863 22695
rect 13863 22661 13872 22695
rect 13820 22652 13872 22661
rect 14096 22652 14148 22704
rect 11520 22584 11572 22636
rect 16028 22627 16080 22636
rect 10784 22516 10836 22568
rect 12716 22516 12768 22568
rect 14372 22559 14424 22568
rect 14372 22525 14381 22559
rect 14381 22525 14415 22559
rect 14415 22525 14424 22559
rect 14372 22516 14424 22525
rect 3240 22380 3292 22432
rect 4068 22380 4120 22432
rect 6184 22380 6236 22432
rect 6920 22423 6972 22432
rect 6920 22389 6929 22423
rect 6929 22389 6963 22423
rect 6963 22389 6972 22423
rect 6920 22380 6972 22389
rect 7288 22380 7340 22432
rect 8760 22423 8812 22432
rect 8760 22389 8769 22423
rect 8769 22389 8803 22423
rect 8803 22389 8812 22423
rect 8760 22380 8812 22389
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 12348 22448 12400 22500
rect 16028 22593 16037 22627
rect 16037 22593 16071 22627
rect 16071 22593 16080 22627
rect 16028 22584 16080 22593
rect 21548 22584 21600 22636
rect 23480 22584 23532 22636
rect 16580 22516 16632 22568
rect 17592 22516 17644 22568
rect 37832 22584 37884 22636
rect 38200 22491 38252 22500
rect 9864 22380 9916 22432
rect 9956 22380 10008 22432
rect 10508 22380 10560 22432
rect 12900 22380 12952 22432
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 15200 22380 15252 22432
rect 17960 22380 18012 22432
rect 38016 22380 38068 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3240 22176 3292 22228
rect 2504 22108 2556 22160
rect 4804 22108 4856 22160
rect 8392 22108 8444 22160
rect 9864 22176 9916 22228
rect 15016 22176 15068 22228
rect 15384 22176 15436 22228
rect 15752 22176 15804 22228
rect 15292 22108 15344 22160
rect 16764 22108 16816 22160
rect 3240 22040 3292 22092
rect 3608 22040 3660 22092
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 3976 21972 4028 22024
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 4620 21972 4672 22024
rect 5080 21972 5132 22024
rect 2964 21947 3016 21956
rect 2964 21913 2973 21947
rect 2973 21913 3007 21947
rect 3007 21913 3016 21947
rect 2964 21904 3016 21913
rect 4436 21904 4488 21956
rect 3240 21836 3292 21888
rect 4160 21836 4212 21888
rect 4712 21836 4764 21888
rect 5724 21904 5776 21956
rect 5908 21836 5960 21888
rect 6552 21972 6604 22024
rect 7012 21904 7064 21956
rect 7656 21972 7708 22024
rect 8116 21972 8168 22024
rect 10048 22040 10100 22092
rect 11796 22040 11848 22092
rect 11888 22040 11940 22092
rect 15108 22083 15160 22092
rect 12440 22015 12492 22024
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12900 22015 12952 22024
rect 12440 21972 12492 21981
rect 12900 21981 12909 22015
rect 12909 21981 12943 22015
rect 12943 21981 12952 22015
rect 12900 21972 12952 21981
rect 13268 21972 13320 22024
rect 15108 22049 15117 22083
rect 15117 22049 15151 22083
rect 15151 22049 15160 22083
rect 15108 22040 15160 22049
rect 15936 22083 15988 22092
rect 15936 22049 15945 22083
rect 15945 22049 15979 22083
rect 15979 22049 15988 22083
rect 15936 22040 15988 22049
rect 17040 22083 17092 22092
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 20260 22176 20312 22228
rect 37832 22219 37884 22228
rect 37832 22185 37841 22219
rect 37841 22185 37875 22219
rect 37875 22185 37884 22219
rect 37832 22176 37884 22185
rect 20168 22108 20220 22160
rect 20352 22108 20404 22160
rect 23112 22040 23164 22092
rect 29000 22040 29052 22092
rect 38016 22015 38068 22024
rect 38016 21981 38025 22015
rect 38025 21981 38059 22015
rect 38059 21981 38068 22015
rect 38016 21972 38068 21981
rect 9220 21947 9272 21956
rect 9220 21913 9229 21947
rect 9229 21913 9263 21947
rect 9263 21913 9272 21947
rect 9220 21904 9272 21913
rect 9312 21947 9364 21956
rect 9312 21913 9321 21947
rect 9321 21913 9355 21947
rect 9355 21913 9364 21947
rect 10784 21947 10836 21956
rect 9312 21904 9364 21913
rect 10784 21913 10793 21947
rect 10793 21913 10827 21947
rect 10827 21913 10836 21947
rect 10784 21904 10836 21913
rect 10876 21947 10928 21956
rect 10876 21913 10885 21947
rect 10885 21913 10919 21947
rect 10919 21913 10928 21947
rect 11428 21947 11480 21956
rect 10876 21904 10928 21913
rect 11428 21913 11437 21947
rect 11437 21913 11471 21947
rect 11471 21913 11480 21947
rect 11428 21904 11480 21913
rect 14556 21904 14608 21956
rect 15200 21947 15252 21956
rect 15200 21913 15209 21947
rect 15209 21913 15243 21947
rect 15243 21913 15252 21947
rect 15200 21904 15252 21913
rect 6552 21836 6604 21888
rect 7564 21836 7616 21888
rect 8300 21836 8352 21888
rect 11888 21836 11940 21888
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 14280 21836 14332 21888
rect 14464 21879 14516 21888
rect 14464 21845 14473 21879
rect 14473 21845 14507 21879
rect 14507 21845 14516 21879
rect 14464 21836 14516 21845
rect 19156 21904 19208 21956
rect 20536 21904 20588 21956
rect 25412 21947 25464 21956
rect 25412 21913 25421 21947
rect 25421 21913 25455 21947
rect 25455 21913 25464 21947
rect 25412 21904 25464 21913
rect 19432 21836 19484 21888
rect 21732 21879 21784 21888
rect 21732 21845 21741 21879
rect 21741 21845 21775 21879
rect 21775 21845 21784 21879
rect 21732 21836 21784 21845
rect 22560 21836 22612 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3240 21632 3292 21684
rect 3976 21632 4028 21684
rect 1860 21607 1912 21616
rect 1860 21573 1869 21607
rect 1869 21573 1903 21607
rect 1903 21573 1912 21607
rect 1860 21564 1912 21573
rect 4160 21564 4212 21616
rect 4896 21632 4948 21684
rect 5080 21632 5132 21684
rect 7196 21607 7248 21616
rect 7196 21573 7205 21607
rect 7205 21573 7239 21607
rect 7239 21573 7248 21607
rect 7196 21564 7248 21573
rect 7380 21564 7432 21616
rect 3608 21428 3660 21480
rect 3792 21471 3844 21480
rect 3792 21437 3801 21471
rect 3801 21437 3835 21471
rect 3835 21437 3844 21471
rect 3792 21428 3844 21437
rect 6828 21496 6880 21548
rect 11060 21632 11112 21684
rect 11428 21632 11480 21684
rect 9772 21564 9824 21616
rect 9864 21564 9916 21616
rect 11612 21564 11664 21616
rect 12256 21564 12308 21616
rect 14464 21564 14516 21616
rect 17132 21564 17184 21616
rect 19156 21607 19208 21616
rect 19156 21573 19165 21607
rect 19165 21573 19199 21607
rect 19199 21573 19208 21607
rect 19156 21564 19208 21573
rect 19984 21564 20036 21616
rect 25412 21632 25464 21684
rect 32312 21675 32364 21684
rect 32312 21641 32321 21675
rect 32321 21641 32355 21675
rect 32355 21641 32364 21675
rect 32312 21632 32364 21641
rect 26240 21564 26292 21616
rect 8852 21428 8904 21480
rect 8944 21428 8996 21480
rect 10600 21496 10652 21548
rect 14188 21496 14240 21548
rect 14924 21496 14976 21548
rect 4712 21360 4764 21412
rect 7288 21360 7340 21412
rect 11152 21428 11204 21480
rect 11888 21428 11940 21480
rect 12716 21428 12768 21480
rect 13268 21471 13320 21480
rect 13268 21437 13277 21471
rect 13277 21437 13311 21471
rect 13311 21437 13320 21471
rect 13268 21428 13320 21437
rect 16120 21428 16172 21480
rect 18328 21428 18380 21480
rect 18604 21496 18656 21548
rect 21732 21496 21784 21548
rect 22192 21539 22244 21548
rect 22192 21505 22201 21539
rect 22201 21505 22235 21539
rect 22235 21505 22244 21539
rect 22192 21496 22244 21505
rect 19800 21471 19852 21480
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 9312 21360 9364 21412
rect 4528 21292 4580 21344
rect 6276 21292 6328 21344
rect 9496 21292 9548 21344
rect 10876 21292 10928 21344
rect 12164 21292 12216 21344
rect 12992 21360 13044 21412
rect 13636 21360 13688 21412
rect 14372 21292 14424 21344
rect 15476 21292 15528 21344
rect 16856 21292 16908 21344
rect 18604 21292 18656 21344
rect 20352 21403 20404 21412
rect 20352 21369 20361 21403
rect 20361 21369 20395 21403
rect 20395 21369 20404 21403
rect 23388 21496 23440 21548
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25136 21496 25188 21505
rect 30472 21496 30524 21548
rect 38016 21539 38068 21548
rect 38016 21505 38025 21539
rect 38025 21505 38059 21539
rect 38059 21505 38068 21539
rect 38016 21496 38068 21505
rect 23112 21471 23164 21480
rect 23112 21437 23121 21471
rect 23121 21437 23155 21471
rect 23155 21437 23164 21471
rect 23112 21428 23164 21437
rect 23664 21428 23716 21480
rect 20352 21360 20404 21369
rect 22376 21335 22428 21344
rect 22376 21301 22385 21335
rect 22385 21301 22419 21335
rect 22419 21301 22428 21335
rect 22376 21292 22428 21301
rect 26332 21360 26384 21412
rect 26516 21403 26568 21412
rect 26516 21369 26525 21403
rect 26525 21369 26559 21403
rect 26559 21369 26568 21403
rect 26516 21360 26568 21369
rect 24400 21292 24452 21344
rect 32404 21360 32456 21412
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1860 21088 1912 21140
rect 2136 21088 2188 21140
rect 2780 21020 2832 21072
rect 3240 21088 3292 21140
rect 4712 21020 4764 21072
rect 7472 21020 7524 21072
rect 8944 21088 8996 21140
rect 9312 21088 9364 21140
rect 9588 21088 9640 21140
rect 11520 21088 11572 21140
rect 16120 21131 16172 21140
rect 9956 21020 10008 21072
rect 6184 20952 6236 21004
rect 8668 20952 8720 21004
rect 8392 20884 8444 20936
rect 9772 20952 9824 21004
rect 11336 21020 11388 21072
rect 12624 21020 12676 21072
rect 12900 21020 12952 21072
rect 13268 21020 13320 21072
rect 14096 21020 14148 21072
rect 14372 21020 14424 21072
rect 15844 21020 15896 21072
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 13176 20952 13228 21004
rect 13636 20952 13688 21004
rect 14648 20995 14700 21004
rect 14648 20961 14657 20995
rect 14657 20961 14691 20995
rect 14691 20961 14700 20995
rect 14648 20952 14700 20961
rect 15016 20952 15068 21004
rect 16120 21097 16129 21131
rect 16129 21097 16163 21131
rect 16163 21097 16172 21131
rect 16120 21088 16172 21097
rect 16212 21088 16264 21140
rect 20536 21131 20588 21140
rect 16028 21020 16080 21072
rect 20536 21097 20545 21131
rect 20545 21097 20579 21131
rect 20579 21097 20588 21131
rect 20536 21088 20588 21097
rect 26240 21131 26292 21140
rect 2320 20859 2372 20868
rect 2320 20825 2329 20859
rect 2329 20825 2363 20859
rect 2363 20825 2372 20859
rect 2320 20816 2372 20825
rect 4528 20816 4580 20868
rect 4804 20859 4856 20868
rect 4804 20825 4813 20859
rect 4813 20825 4847 20859
rect 4847 20825 4856 20859
rect 5908 20859 5960 20868
rect 4804 20816 4856 20825
rect 5908 20825 5917 20859
rect 5917 20825 5951 20859
rect 5951 20825 5960 20859
rect 5908 20816 5960 20825
rect 6000 20859 6052 20868
rect 6000 20825 6009 20859
rect 6009 20825 6043 20859
rect 6043 20825 6052 20859
rect 6000 20816 6052 20825
rect 7288 20816 7340 20868
rect 7564 20859 7616 20868
rect 7564 20825 7573 20859
rect 7573 20825 7607 20859
rect 7607 20825 7616 20859
rect 7564 20816 7616 20825
rect 8300 20816 8352 20868
rect 9220 20816 9272 20868
rect 11152 20884 11204 20936
rect 4896 20748 4948 20800
rect 6552 20748 6604 20800
rect 9864 20816 9916 20868
rect 9680 20748 9732 20800
rect 13636 20816 13688 20868
rect 14556 20816 14608 20868
rect 14740 20816 14792 20868
rect 15200 20884 15252 20936
rect 16948 20952 17000 21004
rect 17224 20995 17276 21004
rect 17224 20961 17233 20995
rect 17233 20961 17267 20995
rect 17267 20961 17276 20995
rect 17224 20952 17276 20961
rect 17408 20952 17460 21004
rect 23756 21020 23808 21072
rect 24124 21020 24176 21072
rect 26240 21097 26249 21131
rect 26249 21097 26283 21131
rect 26283 21097 26292 21131
rect 26240 21088 26292 21097
rect 26332 21088 26384 21140
rect 36084 21088 36136 21140
rect 21732 20952 21784 21004
rect 16212 20884 16264 20936
rect 15936 20816 15988 20868
rect 18420 20884 18472 20936
rect 29920 20952 29972 21004
rect 15200 20748 15252 20800
rect 15384 20748 15436 20800
rect 15752 20748 15804 20800
rect 22376 20816 22428 20868
rect 23848 20816 23900 20868
rect 37188 20884 37240 20936
rect 37832 20884 37884 20936
rect 18144 20748 18196 20800
rect 24860 20791 24912 20800
rect 24860 20757 24869 20791
rect 24869 20757 24903 20791
rect 24903 20757 24912 20791
rect 24860 20748 24912 20757
rect 26792 20791 26844 20800
rect 26792 20757 26801 20791
rect 26801 20757 26835 20791
rect 26835 20757 26844 20791
rect 26792 20748 26844 20757
rect 29920 20748 29972 20800
rect 37740 20748 37792 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1308 20544 1360 20596
rect 2044 20544 2096 20596
rect 1676 20519 1728 20528
rect 1676 20485 1685 20519
rect 1685 20485 1719 20519
rect 1719 20485 1728 20519
rect 1676 20476 1728 20485
rect 1952 20476 2004 20528
rect 2596 20476 2648 20528
rect 4436 20544 4488 20596
rect 4988 20544 5040 20596
rect 3976 20476 4028 20528
rect 7932 20544 7984 20596
rect 8852 20544 8904 20596
rect 6644 20519 6696 20528
rect 6644 20485 6653 20519
rect 6653 20485 6687 20519
rect 6687 20485 6696 20519
rect 6644 20476 6696 20485
rect 7104 20476 7156 20528
rect 8760 20476 8812 20528
rect 6000 20408 6052 20460
rect 3332 20340 3384 20392
rect 5908 20340 5960 20392
rect 6920 20383 6972 20392
rect 6920 20349 6929 20383
rect 6929 20349 6963 20383
rect 6963 20349 6972 20383
rect 6920 20340 6972 20349
rect 9036 20340 9088 20392
rect 9772 20383 9824 20392
rect 4712 20272 4764 20324
rect 6184 20272 6236 20324
rect 6644 20272 6696 20324
rect 9772 20349 9781 20383
rect 9781 20349 9815 20383
rect 9815 20349 9824 20383
rect 9772 20340 9824 20349
rect 10508 20519 10560 20528
rect 10508 20485 10517 20519
rect 10517 20485 10551 20519
rect 10551 20485 10560 20519
rect 10508 20476 10560 20485
rect 11244 20544 11296 20596
rect 12532 20544 12584 20596
rect 10876 20476 10928 20528
rect 13636 20544 13688 20596
rect 13176 20476 13228 20528
rect 13544 20476 13596 20528
rect 15476 20519 15528 20528
rect 15476 20485 15485 20519
rect 15485 20485 15519 20519
rect 15519 20485 15528 20519
rect 15476 20476 15528 20485
rect 15108 20408 15160 20460
rect 12624 20340 12676 20392
rect 15660 20383 15712 20392
rect 6736 20204 6788 20256
rect 7012 20204 7064 20256
rect 8300 20204 8352 20256
rect 9128 20204 9180 20256
rect 9496 20272 9548 20324
rect 10876 20204 10928 20256
rect 12900 20272 12952 20324
rect 13452 20272 13504 20324
rect 15660 20349 15669 20383
rect 15669 20349 15703 20383
rect 15703 20349 15712 20383
rect 15660 20340 15712 20349
rect 22376 20544 22428 20596
rect 23664 20587 23716 20596
rect 23664 20553 23673 20587
rect 23673 20553 23707 20587
rect 23707 20553 23716 20587
rect 23664 20544 23716 20553
rect 23848 20544 23900 20596
rect 17224 20476 17276 20528
rect 26700 20544 26752 20596
rect 25780 20519 25832 20528
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 17960 20408 18012 20460
rect 25780 20485 25789 20519
rect 25789 20485 25823 20519
rect 25823 20485 25832 20519
rect 25780 20476 25832 20485
rect 23572 20451 23624 20460
rect 17868 20340 17920 20392
rect 23572 20417 23581 20451
rect 23581 20417 23615 20451
rect 23615 20417 23624 20451
rect 23572 20408 23624 20417
rect 24400 20451 24452 20460
rect 24400 20417 24409 20451
rect 24409 20417 24443 20451
rect 24443 20417 24452 20451
rect 24400 20408 24452 20417
rect 19064 20272 19116 20324
rect 24860 20340 24912 20392
rect 26516 20340 26568 20392
rect 26976 20340 27028 20392
rect 19524 20272 19576 20324
rect 22560 20272 22612 20324
rect 17316 20204 17368 20256
rect 18880 20204 18932 20256
rect 26884 20204 26936 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4804 20000 4856 20052
rect 6920 19932 6972 19984
rect 9496 19932 9548 19984
rect 4712 19864 4764 19916
rect 4804 19864 4856 19916
rect 6184 19864 6236 19916
rect 8392 19864 8444 19916
rect 10876 20000 10928 20052
rect 15384 20000 15436 20052
rect 16396 20043 16448 20052
rect 16396 20009 16405 20043
rect 16405 20009 16439 20043
rect 16439 20009 16448 20043
rect 16396 20000 16448 20009
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 18328 20000 18380 20052
rect 25780 20043 25832 20052
rect 13176 19932 13228 19984
rect 13820 19932 13872 19984
rect 17132 19932 17184 19984
rect 21640 19932 21692 19984
rect 9772 19864 9824 19916
rect 12072 19907 12124 19916
rect 12072 19873 12081 19907
rect 12081 19873 12115 19907
rect 12115 19873 12124 19907
rect 12072 19864 12124 19873
rect 13544 19907 13596 19916
rect 13544 19873 13553 19907
rect 13553 19873 13587 19907
rect 13587 19873 13596 19907
rect 13544 19864 13596 19873
rect 16672 19864 16724 19916
rect 17316 19864 17368 19916
rect 1860 19796 1912 19848
rect 4344 19839 4396 19848
rect 4344 19805 4353 19839
rect 4353 19805 4387 19839
rect 4387 19805 4396 19839
rect 4344 19796 4396 19805
rect 6552 19796 6604 19848
rect 15752 19796 15804 19848
rect 17500 19796 17552 19848
rect 18604 19796 18656 19848
rect 19524 19796 19576 19848
rect 25780 20009 25789 20043
rect 25789 20009 25823 20043
rect 25823 20009 25832 20043
rect 25780 20000 25832 20009
rect 2504 19771 2556 19780
rect 2504 19737 2513 19771
rect 2513 19737 2547 19771
rect 2547 19737 2556 19771
rect 2504 19728 2556 19737
rect 5172 19771 5224 19780
rect 5172 19737 5181 19771
rect 5181 19737 5215 19771
rect 5215 19737 5224 19771
rect 5172 19728 5224 19737
rect 6184 19728 6236 19780
rect 7012 19771 7064 19780
rect 7012 19737 7021 19771
rect 7021 19737 7055 19771
rect 7055 19737 7064 19771
rect 7012 19728 7064 19737
rect 3700 19660 3752 19712
rect 4712 19660 4764 19712
rect 7656 19771 7708 19780
rect 7656 19737 7665 19771
rect 7665 19737 7699 19771
rect 7699 19737 7708 19771
rect 7656 19728 7708 19737
rect 8944 19660 8996 19712
rect 9404 19771 9456 19780
rect 9404 19737 9413 19771
rect 9413 19737 9447 19771
rect 9447 19737 9456 19771
rect 9404 19728 9456 19737
rect 10140 19728 10192 19780
rect 11520 19771 11572 19780
rect 11520 19737 11529 19771
rect 11529 19737 11563 19771
rect 11563 19737 11572 19771
rect 11520 19728 11572 19737
rect 12164 19771 12216 19780
rect 12164 19737 12173 19771
rect 12173 19737 12207 19771
rect 12207 19737 12216 19771
rect 12164 19728 12216 19737
rect 13176 19728 13228 19780
rect 14464 19771 14516 19780
rect 14464 19737 14473 19771
rect 14473 19737 14507 19771
rect 14507 19737 14516 19771
rect 15384 19771 15436 19780
rect 14464 19728 14516 19737
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 12716 19660 12768 19712
rect 14188 19660 14240 19712
rect 16672 19660 16724 19712
rect 18144 19728 18196 19780
rect 20352 19728 20404 19780
rect 21456 19771 21508 19780
rect 21456 19737 21465 19771
rect 21465 19737 21499 19771
rect 21499 19737 21508 19771
rect 21456 19728 21508 19737
rect 21640 19728 21692 19780
rect 25504 19932 25556 19984
rect 23388 19907 23440 19916
rect 23388 19873 23397 19907
rect 23397 19873 23431 19907
rect 23431 19873 23440 19907
rect 23388 19864 23440 19873
rect 24032 19907 24084 19916
rect 24032 19873 24041 19907
rect 24041 19873 24075 19907
rect 24075 19873 24084 19907
rect 24032 19864 24084 19873
rect 26884 19864 26936 19916
rect 35532 19864 35584 19916
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 26792 19796 26844 19848
rect 26976 19796 27028 19848
rect 23940 19660 23992 19712
rect 24952 19660 25004 19712
rect 34428 19660 34480 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3700 19456 3752 19508
rect 2136 19388 2188 19440
rect 2596 19388 2648 19440
rect 5264 19388 5316 19440
rect 7288 19388 7340 19440
rect 9956 19388 10008 19440
rect 10968 19456 11020 19508
rect 14924 19456 14976 19508
rect 15108 19456 15160 19508
rect 21456 19456 21508 19508
rect 23940 19499 23992 19508
rect 14188 19431 14240 19440
rect 14188 19397 14197 19431
rect 14197 19397 14231 19431
rect 14231 19397 14240 19431
rect 14188 19388 14240 19397
rect 16580 19388 16632 19440
rect 18144 19388 18196 19440
rect 18328 19388 18380 19440
rect 18880 19431 18932 19440
rect 18880 19397 18889 19431
rect 18889 19397 18923 19431
rect 18923 19397 18932 19431
rect 18880 19388 18932 19397
rect 20260 19388 20312 19440
rect 20628 19388 20680 19440
rect 23940 19465 23949 19499
rect 23949 19465 23983 19499
rect 23983 19465 23992 19499
rect 23940 19456 23992 19465
rect 24952 19431 25004 19440
rect 3240 19363 3292 19372
rect 3240 19329 3249 19363
rect 3249 19329 3283 19363
rect 3283 19329 3292 19363
rect 3240 19320 3292 19329
rect 3976 19363 4028 19372
rect 3976 19329 3985 19363
rect 3985 19329 4019 19363
rect 4019 19329 4028 19363
rect 3976 19320 4028 19329
rect 4712 19252 4764 19304
rect 4988 19252 5040 19304
rect 5264 19184 5316 19236
rect 5724 19295 5776 19304
rect 5724 19261 5733 19295
rect 5733 19261 5767 19295
rect 5767 19261 5776 19295
rect 5724 19252 5776 19261
rect 6920 19252 6972 19304
rect 10232 19252 10284 19304
rect 11428 19320 11480 19372
rect 12624 19320 12676 19372
rect 15108 19320 15160 19372
rect 15660 19363 15712 19372
rect 11060 19295 11112 19304
rect 11060 19261 11069 19295
rect 11069 19261 11103 19295
rect 11103 19261 11112 19295
rect 11060 19252 11112 19261
rect 3332 19159 3384 19168
rect 3332 19125 3341 19159
rect 3341 19125 3375 19159
rect 3375 19125 3384 19159
rect 3332 19116 3384 19125
rect 10968 19184 11020 19236
rect 12900 19252 12952 19304
rect 12992 19252 13044 19304
rect 13544 19252 13596 19304
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 19340 19320 19392 19372
rect 22192 19363 22244 19372
rect 17868 19295 17920 19304
rect 13176 19184 13228 19236
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 15292 19184 15344 19236
rect 15844 19184 15896 19236
rect 21916 19184 21968 19236
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 24952 19397 24961 19431
rect 24961 19397 24995 19431
rect 24995 19397 25004 19431
rect 24952 19388 25004 19397
rect 25504 19431 25556 19440
rect 25504 19397 25513 19431
rect 25513 19397 25547 19431
rect 25547 19397 25556 19431
rect 25504 19388 25556 19397
rect 38292 19363 38344 19372
rect 38292 19329 38301 19363
rect 38301 19329 38335 19363
rect 38335 19329 38344 19363
rect 38292 19320 38344 19329
rect 24860 19295 24912 19304
rect 24860 19261 24869 19295
rect 24869 19261 24903 19295
rect 24903 19261 24912 19295
rect 24860 19252 24912 19261
rect 24952 19252 25004 19304
rect 8024 19116 8076 19168
rect 8392 19116 8444 19168
rect 9312 19116 9364 19168
rect 12532 19116 12584 19168
rect 13728 19116 13780 19168
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 23388 19116 23440 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3424 18912 3476 18964
rect 8576 18955 8628 18964
rect 8576 18921 8585 18955
rect 8585 18921 8619 18955
rect 8619 18921 8628 18955
rect 8576 18912 8628 18921
rect 8668 18912 8720 18964
rect 9956 18912 10008 18964
rect 15568 18955 15620 18964
rect 15568 18921 15577 18955
rect 15577 18921 15611 18955
rect 15611 18921 15620 18955
rect 15568 18912 15620 18921
rect 17224 18955 17276 18964
rect 17224 18921 17233 18955
rect 17233 18921 17267 18955
rect 17267 18921 17276 18955
rect 17224 18912 17276 18921
rect 19432 18912 19484 18964
rect 22836 18912 22888 18964
rect 8944 18844 8996 18896
rect 9036 18844 9088 18896
rect 3332 18776 3384 18828
rect 14556 18776 14608 18828
rect 16764 18776 16816 18828
rect 1584 18751 1636 18760
rect 1584 18717 1593 18751
rect 1593 18717 1627 18751
rect 1627 18717 1636 18751
rect 1584 18708 1636 18717
rect 3976 18708 4028 18760
rect 6552 18708 6604 18760
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 3148 18640 3200 18692
rect 7104 18683 7156 18692
rect 7104 18649 7113 18683
rect 7113 18649 7147 18683
rect 7147 18649 7156 18683
rect 7104 18640 7156 18649
rect 7380 18640 7432 18692
rect 3792 18572 3844 18624
rect 6000 18572 6052 18624
rect 7472 18572 7524 18624
rect 10048 18708 10100 18760
rect 10508 18708 10560 18760
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 12440 18708 12492 18760
rect 14096 18708 14148 18760
rect 16028 18708 16080 18760
rect 16396 18708 16448 18760
rect 24032 18776 24084 18828
rect 24952 18819 25004 18828
rect 24952 18785 24961 18819
rect 24961 18785 24995 18819
rect 24995 18785 25004 18819
rect 24952 18776 25004 18785
rect 19984 18708 20036 18760
rect 20260 18751 20312 18760
rect 20260 18717 20269 18751
rect 20269 18717 20303 18751
rect 20303 18717 20312 18751
rect 20260 18708 20312 18717
rect 25044 18708 25096 18760
rect 9588 18640 9640 18692
rect 10692 18683 10744 18692
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 10048 18615 10100 18624
rect 9404 18572 9456 18581
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 10692 18649 10701 18683
rect 10701 18649 10735 18683
rect 10735 18649 10744 18683
rect 10692 18640 10744 18649
rect 10784 18683 10836 18692
rect 10784 18649 10793 18683
rect 10793 18649 10827 18683
rect 10827 18649 10836 18683
rect 11704 18683 11756 18692
rect 10784 18640 10836 18649
rect 11704 18649 11713 18683
rect 11713 18649 11747 18683
rect 11747 18649 11756 18683
rect 11704 18640 11756 18649
rect 12348 18640 12400 18692
rect 14188 18640 14240 18692
rect 11980 18572 12032 18624
rect 14280 18572 14332 18624
rect 14556 18640 14608 18692
rect 18420 18640 18472 18692
rect 22836 18640 22888 18692
rect 23204 18640 23256 18692
rect 38016 18844 38068 18896
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 20536 18572 20588 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2780 18368 2832 18420
rect 3332 18411 3384 18420
rect 3332 18377 3341 18411
rect 3341 18377 3375 18411
rect 3375 18377 3384 18411
rect 3332 18368 3384 18377
rect 4068 18368 4120 18420
rect 4620 18300 4672 18352
rect 5448 18232 5500 18284
rect 6828 18368 6880 18420
rect 6736 18300 6788 18352
rect 9312 18343 9364 18352
rect 9312 18309 9321 18343
rect 9321 18309 9355 18343
rect 9355 18309 9364 18343
rect 9312 18300 9364 18309
rect 10048 18300 10100 18352
rect 11060 18300 11112 18352
rect 11520 18300 11572 18352
rect 11704 18368 11756 18420
rect 12992 18368 13044 18420
rect 11888 18300 11940 18352
rect 12072 18300 12124 18352
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 3424 18164 3476 18216
rect 5724 18164 5776 18216
rect 6092 18164 6144 18216
rect 2872 18096 2924 18148
rect 6920 18164 6972 18216
rect 8944 18164 8996 18216
rect 9864 18164 9916 18216
rect 9956 18164 10008 18216
rect 10784 18232 10836 18284
rect 14924 18368 14976 18420
rect 15016 18368 15068 18420
rect 21180 18368 21232 18420
rect 23204 18411 23256 18420
rect 23204 18377 23213 18411
rect 23213 18377 23247 18411
rect 23247 18377 23256 18411
rect 23204 18368 23256 18377
rect 24400 18368 24452 18420
rect 25044 18411 25096 18420
rect 25044 18377 25053 18411
rect 25053 18377 25087 18411
rect 25087 18377 25096 18411
rect 25044 18368 25096 18377
rect 13452 18300 13504 18352
rect 14280 18300 14332 18352
rect 15016 18232 15068 18284
rect 18236 18300 18288 18352
rect 20628 18300 20680 18352
rect 17960 18232 18012 18284
rect 23388 18275 23440 18284
rect 23388 18241 23397 18275
rect 23397 18241 23431 18275
rect 23431 18241 23440 18275
rect 23388 18232 23440 18241
rect 24032 18275 24084 18284
rect 24032 18241 24041 18275
rect 24041 18241 24075 18275
rect 24075 18241 24084 18275
rect 24032 18232 24084 18241
rect 25688 18275 25740 18284
rect 10692 18164 10744 18216
rect 11520 18164 11572 18216
rect 14464 18164 14516 18216
rect 16948 18164 17000 18216
rect 19248 18164 19300 18216
rect 21916 18164 21968 18216
rect 23572 18164 23624 18216
rect 25688 18241 25697 18275
rect 25697 18241 25731 18275
rect 25731 18241 25740 18275
rect 25688 18232 25740 18241
rect 34428 18232 34480 18284
rect 35440 18232 35492 18284
rect 15016 18096 15068 18148
rect 19984 18096 20036 18148
rect 10692 18028 10744 18080
rect 10876 18028 10928 18080
rect 11244 18028 11296 18080
rect 13452 18071 13504 18080
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 13544 18028 13596 18080
rect 15936 18028 15988 18080
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 18328 18028 18380 18080
rect 25780 18071 25832 18080
rect 25780 18037 25789 18071
rect 25789 18037 25823 18071
rect 25823 18037 25832 18071
rect 25780 18028 25832 18037
rect 38016 18028 38068 18080
rect 38200 18071 38252 18080
rect 38200 18037 38209 18071
rect 38209 18037 38243 18071
rect 38243 18037 38252 18071
rect 38200 18028 38252 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3976 17824 4028 17876
rect 4068 17824 4120 17876
rect 3056 17756 3108 17808
rect 3792 17756 3844 17808
rect 1676 17731 1728 17740
rect 1676 17697 1685 17731
rect 1685 17697 1719 17731
rect 1719 17697 1728 17731
rect 5448 17756 5500 17808
rect 10784 17824 10836 17876
rect 12072 17824 12124 17876
rect 12256 17824 12308 17876
rect 15844 17824 15896 17876
rect 16580 17824 16632 17876
rect 18788 17824 18840 17876
rect 1676 17688 1728 17697
rect 4712 17688 4764 17740
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 8944 17688 8996 17740
rect 11520 17688 11572 17740
rect 12256 17688 12308 17740
rect 12348 17688 12400 17740
rect 15016 17688 15068 17740
rect 1952 17595 2004 17604
rect 1952 17561 1961 17595
rect 1961 17561 1995 17595
rect 1995 17561 2004 17595
rect 1952 17552 2004 17561
rect 4252 17552 4304 17604
rect 5080 17552 5132 17604
rect 4988 17484 5040 17536
rect 5908 17484 5960 17536
rect 9312 17552 9364 17604
rect 9128 17484 9180 17536
rect 10968 17552 11020 17604
rect 10876 17484 10928 17536
rect 15292 17620 15344 17672
rect 22652 17756 22704 17808
rect 20352 17688 20404 17740
rect 21272 17688 21324 17740
rect 11888 17595 11940 17604
rect 11888 17561 11897 17595
rect 11897 17561 11931 17595
rect 11931 17561 11940 17595
rect 11888 17552 11940 17561
rect 13176 17552 13228 17604
rect 14188 17552 14240 17604
rect 14464 17595 14516 17604
rect 14464 17561 14473 17595
rect 14473 17561 14507 17595
rect 14507 17561 14516 17595
rect 15384 17595 15436 17604
rect 14464 17552 14516 17561
rect 15384 17561 15393 17595
rect 15393 17561 15427 17595
rect 15427 17561 15436 17595
rect 15384 17552 15436 17561
rect 17500 17552 17552 17604
rect 13820 17484 13872 17536
rect 14832 17484 14884 17536
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 17224 17527 17276 17536
rect 17224 17493 17233 17527
rect 17233 17493 17267 17527
rect 17267 17493 17276 17527
rect 17224 17484 17276 17493
rect 20076 17552 20128 17604
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2596 17280 2648 17332
rect 1860 17255 1912 17264
rect 1860 17221 1869 17255
rect 1869 17221 1903 17255
rect 1903 17221 1912 17255
rect 1860 17212 1912 17221
rect 4068 17212 4120 17264
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 1952 17076 2004 17128
rect 3792 17144 3844 17196
rect 3608 17119 3660 17128
rect 3608 17085 3617 17119
rect 3617 17085 3651 17119
rect 3651 17085 3660 17119
rect 3608 17076 3660 17085
rect 2964 17008 3016 17060
rect 3976 17008 4028 17060
rect 1492 16940 1544 16992
rect 6092 17280 6144 17332
rect 4528 17255 4580 17264
rect 4528 17221 4537 17255
rect 4537 17221 4571 17255
rect 4571 17221 4580 17255
rect 4528 17212 4580 17221
rect 10048 17280 10100 17332
rect 5632 17144 5684 17196
rect 4620 17076 4672 17128
rect 4896 17076 4948 17128
rect 7104 17076 7156 17128
rect 8576 17076 8628 17128
rect 9680 17144 9732 17196
rect 10048 17187 10100 17196
rect 10048 17153 10057 17187
rect 10057 17153 10091 17187
rect 10091 17153 10100 17187
rect 10048 17144 10100 17153
rect 10692 17212 10744 17264
rect 11980 17255 12032 17264
rect 11980 17221 11989 17255
rect 11989 17221 12023 17255
rect 12023 17221 12032 17255
rect 11980 17212 12032 17221
rect 12072 17212 12124 17264
rect 14464 17280 14516 17332
rect 35440 17280 35492 17332
rect 15200 17212 15252 17264
rect 17224 17212 17276 17264
rect 23940 17212 23992 17264
rect 25780 17212 25832 17264
rect 11336 17144 11388 17196
rect 10876 17076 10928 17128
rect 9312 17008 9364 17060
rect 11612 17008 11664 17060
rect 5080 16940 5132 16992
rect 6368 16940 6420 16992
rect 6736 16983 6788 16992
rect 6736 16949 6745 16983
rect 6745 16949 6779 16983
rect 6779 16949 6788 16983
rect 6736 16940 6788 16949
rect 11428 16940 11480 16992
rect 11520 16940 11572 16992
rect 13636 17144 13688 17196
rect 14740 17076 14792 17128
rect 15384 16940 15436 16992
rect 16396 17008 16448 17060
rect 19432 17144 19484 17196
rect 23756 17144 23808 17196
rect 31760 17144 31812 17196
rect 23020 17119 23072 17128
rect 23020 17085 23029 17119
rect 23029 17085 23063 17119
rect 23063 17085 23072 17119
rect 23020 17076 23072 17085
rect 24400 17119 24452 17128
rect 24400 17085 24409 17119
rect 24409 17085 24443 17119
rect 24443 17085 24452 17119
rect 24400 17076 24452 17085
rect 25688 17076 25740 17128
rect 17040 17008 17092 17060
rect 24032 17008 24084 17060
rect 16856 16940 16908 16992
rect 17684 16940 17736 16992
rect 18052 16940 18104 16992
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 20904 16940 20956 16992
rect 26148 16940 26200 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1492 16736 1544 16788
rect 1584 16736 1636 16788
rect 2044 16736 2096 16788
rect 6092 16736 6144 16788
rect 6368 16736 6420 16788
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 4160 16668 4212 16720
rect 4896 16668 4948 16720
rect 9312 16779 9364 16788
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 9956 16736 10008 16788
rect 11796 16736 11848 16788
rect 3608 16600 3660 16652
rect 3884 16532 3936 16584
rect 4620 16600 4672 16652
rect 7104 16600 7156 16652
rect 9588 16668 9640 16720
rect 11060 16668 11112 16720
rect 12716 16668 12768 16720
rect 12900 16711 12952 16720
rect 12900 16677 12909 16711
rect 12909 16677 12943 16711
rect 12943 16677 12952 16711
rect 12900 16668 12952 16677
rect 13176 16736 13228 16788
rect 15844 16736 15896 16788
rect 16120 16736 16172 16788
rect 19340 16736 19392 16788
rect 17040 16668 17092 16720
rect 37924 16736 37976 16788
rect 5080 16532 5132 16584
rect 8576 16532 8628 16584
rect 9588 16532 9640 16584
rect 11520 16600 11572 16652
rect 11888 16600 11940 16652
rect 12164 16600 12216 16652
rect 12992 16600 13044 16652
rect 13360 16600 13412 16652
rect 10140 16532 10192 16584
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 16764 16600 16816 16652
rect 18328 16643 18380 16652
rect 18328 16609 18337 16643
rect 18337 16609 18371 16643
rect 18371 16609 18380 16643
rect 18328 16600 18380 16609
rect 10508 16532 10560 16541
rect 14096 16532 14148 16584
rect 3976 16507 4028 16516
rect 3976 16473 3985 16507
rect 3985 16473 4019 16507
rect 4019 16473 4028 16507
rect 3976 16464 4028 16473
rect 4252 16464 4304 16516
rect 4712 16507 4764 16516
rect 4712 16473 4721 16507
rect 4721 16473 4755 16507
rect 4755 16473 4764 16507
rect 4712 16464 4764 16473
rect 5632 16464 5684 16516
rect 7656 16507 7708 16516
rect 2872 16396 2924 16448
rect 7656 16473 7665 16507
rect 7665 16473 7699 16507
rect 7699 16473 7708 16507
rect 7656 16464 7708 16473
rect 9680 16464 9732 16516
rect 8024 16396 8076 16448
rect 9588 16396 9640 16448
rect 11152 16464 11204 16516
rect 14832 16464 14884 16516
rect 15016 16507 15068 16516
rect 15016 16473 15025 16507
rect 15025 16473 15059 16507
rect 15059 16473 15068 16507
rect 15016 16464 15068 16473
rect 15568 16532 15620 16584
rect 18604 16532 18656 16584
rect 15844 16464 15896 16516
rect 16764 16507 16816 16516
rect 16764 16473 16773 16507
rect 16773 16473 16807 16507
rect 16807 16473 16816 16507
rect 17684 16507 17736 16516
rect 16764 16464 16816 16473
rect 17684 16473 17693 16507
rect 17693 16473 17727 16507
rect 17727 16473 17736 16507
rect 17684 16464 17736 16473
rect 19984 16532 20036 16584
rect 20812 16575 20864 16584
rect 20812 16541 20821 16575
rect 20821 16541 20855 16575
rect 20855 16541 20864 16575
rect 20812 16532 20864 16541
rect 22192 16532 22244 16584
rect 22928 16532 22980 16584
rect 24032 16600 24084 16652
rect 24860 16600 24912 16652
rect 25504 16600 25556 16652
rect 26148 16643 26200 16652
rect 26148 16609 26157 16643
rect 26157 16609 26191 16643
rect 26191 16609 26200 16643
rect 26148 16600 26200 16609
rect 27712 16600 27764 16652
rect 23940 16575 23992 16584
rect 23940 16541 23949 16575
rect 23949 16541 23983 16575
rect 23983 16541 23992 16575
rect 23940 16532 23992 16541
rect 21456 16464 21508 16516
rect 23388 16464 23440 16516
rect 24768 16507 24820 16516
rect 24768 16473 24777 16507
rect 24777 16473 24811 16507
rect 24811 16473 24820 16507
rect 25688 16507 25740 16516
rect 24768 16464 24820 16473
rect 25688 16473 25697 16507
rect 25697 16473 25731 16507
rect 25731 16473 25740 16507
rect 25688 16464 25740 16473
rect 31760 16532 31812 16584
rect 38016 16575 38068 16584
rect 38016 16541 38025 16575
rect 38025 16541 38059 16575
rect 38059 16541 38068 16575
rect 38016 16532 38068 16541
rect 10876 16396 10928 16448
rect 17960 16396 18012 16448
rect 19984 16439 20036 16448
rect 19984 16405 19993 16439
rect 19993 16405 20027 16439
rect 20027 16405 20036 16439
rect 19984 16396 20036 16405
rect 20260 16396 20312 16448
rect 22008 16396 22060 16448
rect 24400 16396 24452 16448
rect 26792 16439 26844 16448
rect 26792 16405 26801 16439
rect 26801 16405 26835 16439
rect 26835 16405 26844 16439
rect 26792 16396 26844 16405
rect 38200 16439 38252 16448
rect 38200 16405 38209 16439
rect 38209 16405 38243 16439
rect 38243 16405 38252 16439
rect 38200 16396 38252 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3792 16192 3844 16244
rect 6000 16235 6052 16244
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 9588 16192 9640 16244
rect 10784 16192 10836 16244
rect 12900 16192 12952 16244
rect 13268 16192 13320 16244
rect 20812 16235 20864 16244
rect 3332 16124 3384 16176
rect 5816 16124 5868 16176
rect 7656 16124 7708 16176
rect 11336 16124 11388 16176
rect 1676 16056 1728 16108
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 9772 16056 9824 16108
rect 10416 16056 10468 16108
rect 10508 16099 10560 16108
rect 10508 16065 10517 16099
rect 10517 16065 10551 16099
rect 10551 16065 10560 16099
rect 10508 16056 10560 16065
rect 2780 15988 2832 16040
rect 5540 15988 5592 16040
rect 6184 15988 6236 16040
rect 10324 15988 10376 16040
rect 12256 16124 12308 16176
rect 11520 15988 11572 16040
rect 13360 15988 13412 16040
rect 9864 15920 9916 15972
rect 6092 15852 6144 15904
rect 9128 15852 9180 15904
rect 9220 15852 9272 15904
rect 10324 15852 10376 15904
rect 11980 15852 12032 15904
rect 13360 15852 13412 15904
rect 14832 16124 14884 16176
rect 17316 16124 17368 16176
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 24768 16192 24820 16244
rect 27712 16235 27764 16244
rect 27712 16201 27721 16235
rect 27721 16201 27755 16235
rect 27755 16201 27764 16235
rect 27712 16192 27764 16201
rect 22192 16167 22244 16176
rect 22192 16133 22201 16167
rect 22201 16133 22235 16167
rect 22235 16133 22244 16167
rect 22192 16124 22244 16133
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 14740 16056 14792 16108
rect 15568 16056 15620 16108
rect 15844 16056 15896 16108
rect 16304 16056 16356 16108
rect 13820 15988 13872 16040
rect 14556 15920 14608 15972
rect 16580 15988 16632 16040
rect 18972 16056 19024 16108
rect 19432 15988 19484 16040
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 27620 16099 27672 16108
rect 27620 16065 27629 16099
rect 27629 16065 27663 16099
rect 27663 16065 27672 16099
rect 27620 16056 27672 16065
rect 36544 16056 36596 16108
rect 15384 15920 15436 15972
rect 17500 15963 17552 15972
rect 17500 15929 17509 15963
rect 17509 15929 17543 15963
rect 17543 15929 17552 15963
rect 17500 15920 17552 15929
rect 17684 15920 17736 15972
rect 18880 15920 18932 15972
rect 21824 15988 21876 16040
rect 21732 15920 21784 15972
rect 24584 15988 24636 16040
rect 18512 15852 18564 15904
rect 18696 15852 18748 15904
rect 25688 15920 25740 15972
rect 24768 15852 24820 15904
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3608 15648 3660 15700
rect 7196 15648 7248 15700
rect 11796 15691 11848 15700
rect 5540 15580 5592 15632
rect 6092 15580 6144 15632
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 12440 15648 12492 15700
rect 14740 15648 14792 15700
rect 16580 15648 16632 15700
rect 21732 15648 21784 15700
rect 22468 15691 22520 15700
rect 22468 15657 22477 15691
rect 22477 15657 22511 15691
rect 22511 15657 22520 15691
rect 22468 15648 22520 15657
rect 23020 15648 23072 15700
rect 26792 15648 26844 15700
rect 13544 15580 13596 15632
rect 15568 15623 15620 15632
rect 15568 15589 15577 15623
rect 15577 15589 15611 15623
rect 15611 15589 15620 15623
rect 15568 15580 15620 15589
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 3424 15512 3476 15564
rect 4620 15512 4672 15564
rect 6828 15512 6880 15564
rect 10692 15512 10744 15564
rect 11612 15512 11664 15564
rect 12808 15512 12860 15564
rect 13176 15512 13228 15564
rect 5356 15444 5408 15496
rect 1952 15308 2004 15360
rect 2596 15308 2648 15360
rect 4160 15376 4212 15428
rect 6460 15376 6512 15428
rect 6736 15376 6788 15428
rect 6184 15308 6236 15360
rect 7840 15376 7892 15428
rect 12256 15444 12308 15496
rect 12532 15444 12584 15496
rect 18696 15512 18748 15564
rect 6920 15308 6972 15360
rect 7748 15308 7800 15360
rect 8484 15308 8536 15360
rect 9588 15308 9640 15360
rect 10324 15419 10376 15428
rect 10324 15385 10333 15419
rect 10333 15385 10367 15419
rect 10367 15385 10376 15419
rect 10324 15376 10376 15385
rect 11060 15376 11112 15428
rect 12440 15308 12492 15360
rect 12900 15376 12952 15428
rect 15016 15376 15068 15428
rect 15200 15444 15252 15496
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 15292 15376 15344 15428
rect 15844 15376 15896 15428
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17868 15487 17920 15496
rect 17316 15444 17368 15453
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 18420 15444 18472 15496
rect 20812 15580 20864 15632
rect 21548 15580 21600 15632
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 23388 15580 23440 15632
rect 27988 15580 28040 15632
rect 24584 15555 24636 15564
rect 14832 15308 14884 15360
rect 17040 15308 17092 15360
rect 17132 15308 17184 15360
rect 19340 15376 19392 15428
rect 19984 15376 20036 15428
rect 20352 15376 20404 15428
rect 22928 15376 22980 15428
rect 17960 15351 18012 15360
rect 17960 15317 17969 15351
rect 17969 15317 18003 15351
rect 18003 15317 18012 15351
rect 17960 15308 18012 15317
rect 18604 15351 18656 15360
rect 18604 15317 18613 15351
rect 18613 15317 18647 15351
rect 18647 15317 18656 15351
rect 18604 15308 18656 15317
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 21548 15308 21600 15360
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 24768 15555 24820 15564
rect 24768 15521 24777 15555
rect 24777 15521 24811 15555
rect 24811 15521 24820 15555
rect 24768 15512 24820 15521
rect 28816 15308 28868 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 3608 15104 3660 15156
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 4160 15036 4212 15088
rect 8484 15104 8536 15156
rect 9128 15104 9180 15156
rect 4988 15036 5040 15088
rect 7840 15036 7892 15088
rect 2412 14900 2464 14952
rect 2596 14900 2648 14952
rect 7104 14968 7156 15020
rect 7472 14968 7524 15020
rect 9956 15104 10008 15156
rect 10232 15036 10284 15088
rect 12900 15104 12952 15156
rect 13360 15104 13412 15156
rect 17960 15104 18012 15156
rect 18512 15147 18564 15156
rect 18512 15113 18521 15147
rect 18521 15113 18555 15147
rect 18555 15113 18564 15147
rect 18512 15104 18564 15113
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 22192 15104 22244 15156
rect 15016 15036 15068 15088
rect 17040 15079 17092 15088
rect 17040 15045 17049 15079
rect 17049 15045 17083 15079
rect 17083 15045 17092 15079
rect 17040 15036 17092 15045
rect 20904 15036 20956 15088
rect 21824 15036 21876 15088
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 20168 14968 20220 15020
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 23848 14968 23900 15020
rect 26056 14968 26108 15020
rect 28816 15011 28868 15020
rect 28816 14977 28825 15011
rect 28825 14977 28859 15011
rect 28859 14977 28868 15011
rect 28816 14968 28868 14977
rect 37832 14968 37884 15020
rect 3332 14943 3384 14952
rect 3332 14909 3341 14943
rect 3341 14909 3375 14943
rect 3375 14909 3384 14943
rect 3332 14900 3384 14909
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 6828 14900 6880 14952
rect 9956 14900 10008 14952
rect 11520 14900 11572 14952
rect 12072 14900 12124 14952
rect 15568 14900 15620 14952
rect 17592 14943 17644 14952
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 19340 14900 19392 14952
rect 7012 14832 7064 14884
rect 4712 14764 4764 14816
rect 5632 14764 5684 14816
rect 7472 14807 7524 14816
rect 7472 14773 7481 14807
rect 7481 14773 7515 14807
rect 7515 14773 7524 14807
rect 7472 14764 7524 14773
rect 10140 14832 10192 14884
rect 10508 14832 10560 14884
rect 26148 14900 26200 14952
rect 26700 14900 26752 14952
rect 9772 14764 9824 14816
rect 10048 14764 10100 14816
rect 10784 14764 10836 14816
rect 11244 14764 11296 14816
rect 13820 14764 13872 14816
rect 15292 14764 15344 14816
rect 18420 14764 18472 14816
rect 24768 14764 24820 14816
rect 26792 14764 26844 14816
rect 37924 14764 37976 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 7196 14603 7248 14612
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 4804 14492 4856 14544
rect 5448 14492 5500 14544
rect 7196 14569 7205 14603
rect 7205 14569 7239 14603
rect 7239 14569 7248 14603
rect 7196 14560 7248 14569
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 8024 14560 8076 14612
rect 9864 14560 9916 14612
rect 9956 14560 10008 14612
rect 8668 14492 8720 14544
rect 10416 14492 10468 14544
rect 4252 14424 4304 14476
rect 5724 14467 5776 14476
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 6460 14424 6512 14476
rect 4896 14356 4948 14408
rect 5448 14399 5500 14408
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 7564 14356 7616 14408
rect 8024 14356 8076 14408
rect 2596 14220 2648 14272
rect 5632 14220 5684 14272
rect 6736 14288 6788 14340
rect 7196 14220 7248 14272
rect 8392 14220 8444 14272
rect 8852 14356 8904 14408
rect 11520 14424 11572 14476
rect 13912 14492 13964 14544
rect 16764 14560 16816 14612
rect 18236 14560 18288 14612
rect 20628 14603 20680 14612
rect 15108 14492 15160 14544
rect 15200 14424 15252 14476
rect 15476 14467 15528 14476
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 15568 14424 15620 14476
rect 18604 14424 18656 14476
rect 18972 14424 19024 14476
rect 10692 14356 10744 14408
rect 10784 14356 10836 14408
rect 9404 14331 9456 14340
rect 9404 14297 9413 14331
rect 9413 14297 9447 14331
rect 9447 14297 9456 14331
rect 9404 14288 9456 14297
rect 9496 14288 9548 14340
rect 14464 14356 14516 14408
rect 18144 14356 18196 14408
rect 20628 14569 20637 14603
rect 20637 14569 20671 14603
rect 20671 14569 20680 14603
rect 20628 14560 20680 14569
rect 21272 14560 21324 14612
rect 34520 14560 34572 14612
rect 36544 14560 36596 14612
rect 20904 14492 20956 14544
rect 21456 14492 21508 14544
rect 20260 14424 20312 14476
rect 22008 14424 22060 14476
rect 24768 14467 24820 14476
rect 24768 14433 24777 14467
rect 24777 14433 24811 14467
rect 24811 14433 24820 14467
rect 24768 14424 24820 14433
rect 26700 14467 26752 14476
rect 26700 14433 26709 14467
rect 26709 14433 26743 14467
rect 26743 14433 26752 14467
rect 26700 14424 26752 14433
rect 21548 14356 21600 14408
rect 21916 14356 21968 14408
rect 26148 14356 26200 14408
rect 27988 14399 28040 14408
rect 27988 14365 27997 14399
rect 27997 14365 28031 14399
rect 28031 14365 28040 14399
rect 27988 14356 28040 14365
rect 34612 14356 34664 14408
rect 37280 14356 37332 14408
rect 11796 14288 11848 14340
rect 11980 14288 12032 14340
rect 10324 14220 10376 14272
rect 10416 14220 10468 14272
rect 17868 14288 17920 14340
rect 17040 14220 17092 14272
rect 17776 14220 17828 14272
rect 20352 14288 20404 14340
rect 18696 14220 18748 14272
rect 20904 14220 20956 14272
rect 26608 14220 26660 14272
rect 27344 14263 27396 14272
rect 27344 14229 27353 14263
rect 27353 14229 27387 14263
rect 27387 14229 27396 14263
rect 27344 14220 27396 14229
rect 28080 14263 28132 14272
rect 28080 14229 28089 14263
rect 28089 14229 28123 14263
rect 28123 14229 28132 14263
rect 28080 14220 28132 14229
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2780 14016 2832 14068
rect 13452 14059 13504 14068
rect 6460 13948 6512 14000
rect 7380 13948 7432 14000
rect 7472 13948 7524 14000
rect 10048 13948 10100 14000
rect 10416 13991 10468 14000
rect 10416 13957 10425 13991
rect 10425 13957 10459 13991
rect 10459 13957 10468 13991
rect 10416 13948 10468 13957
rect 11060 13991 11112 14000
rect 11060 13957 11069 13991
rect 11069 13957 11103 13991
rect 11103 13957 11112 13991
rect 11060 13948 11112 13957
rect 12440 13948 12492 14000
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 15016 14016 15068 14068
rect 14096 13991 14148 14000
rect 14096 13957 14105 13991
rect 14105 13957 14139 13991
rect 14139 13957 14148 13991
rect 14096 13948 14148 13957
rect 14280 13948 14332 14000
rect 15200 13948 15252 14000
rect 17040 13991 17092 14000
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 4160 13880 4212 13932
rect 7196 13923 7248 13932
rect 2688 13812 2740 13864
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 5264 13812 5316 13864
rect 6276 13812 6328 13864
rect 7196 13889 7205 13923
rect 7205 13889 7239 13923
rect 7239 13889 7248 13923
rect 7196 13880 7248 13889
rect 9496 13880 9548 13932
rect 10508 13880 10560 13932
rect 10784 13880 10836 13932
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 17040 13957 17049 13991
rect 17049 13957 17083 13991
rect 17083 13957 17092 13991
rect 17040 13948 17092 13957
rect 20536 14016 20588 14068
rect 17684 13948 17736 14000
rect 18696 13991 18748 14000
rect 18696 13957 18705 13991
rect 18705 13957 18739 13991
rect 18739 13957 18748 13991
rect 18696 13948 18748 13957
rect 22468 14016 22520 14068
rect 26608 14059 26660 14068
rect 26608 14025 26617 14059
rect 26617 14025 26651 14059
rect 26651 14025 26660 14059
rect 26608 14016 26660 14025
rect 20812 13923 20864 13932
rect 7472 13812 7524 13864
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 6736 13744 6788 13796
rect 9404 13812 9456 13864
rect 10048 13812 10100 13864
rect 11980 13855 12032 13864
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 14648 13812 14700 13864
rect 15476 13812 15528 13864
rect 17500 13812 17552 13864
rect 20812 13889 20821 13923
rect 20821 13889 20855 13923
rect 20855 13889 20864 13923
rect 20812 13880 20864 13889
rect 22376 13880 22428 13932
rect 23572 13923 23624 13932
rect 23572 13889 23581 13923
rect 23581 13889 23615 13923
rect 23615 13889 23624 13923
rect 23572 13880 23624 13889
rect 26792 13948 26844 14000
rect 34796 14016 34848 14068
rect 27344 13923 27396 13932
rect 27344 13889 27353 13923
rect 27353 13889 27387 13923
rect 27387 13889 27396 13923
rect 27344 13880 27396 13889
rect 18788 13812 18840 13864
rect 19708 13855 19760 13864
rect 19708 13821 19717 13855
rect 19717 13821 19751 13855
rect 19751 13821 19760 13855
rect 19708 13812 19760 13821
rect 22100 13812 22152 13864
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 26608 13812 26660 13864
rect 4620 13676 4672 13728
rect 7196 13676 7248 13728
rect 10232 13744 10284 13796
rect 17224 13744 17276 13796
rect 13912 13676 13964 13728
rect 15108 13676 15160 13728
rect 16120 13676 16172 13728
rect 20996 13744 21048 13796
rect 21088 13744 21140 13796
rect 23296 13744 23348 13796
rect 19708 13676 19760 13728
rect 22928 13676 22980 13728
rect 23388 13719 23440 13728
rect 23388 13685 23397 13719
rect 23397 13685 23431 13719
rect 23431 13685 23440 13719
rect 23388 13676 23440 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2964 13472 3016 13524
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 5356 13472 5408 13524
rect 6092 13472 6144 13524
rect 9496 13472 9548 13524
rect 9956 13472 10008 13524
rect 11980 13472 12032 13524
rect 14464 13472 14516 13524
rect 9036 13404 9088 13456
rect 13636 13404 13688 13456
rect 18236 13472 18288 13524
rect 20076 13472 20128 13524
rect 20536 13472 20588 13524
rect 22468 13515 22520 13524
rect 22468 13481 22477 13515
rect 22477 13481 22511 13515
rect 22511 13481 22520 13515
rect 22468 13472 22520 13481
rect 26792 13515 26844 13524
rect 26792 13481 26801 13515
rect 26801 13481 26835 13515
rect 26835 13481 26844 13515
rect 26792 13472 26844 13481
rect 18052 13404 18104 13456
rect 20444 13404 20496 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 4620 13336 4672 13388
rect 6552 13336 6604 13388
rect 8944 13336 8996 13388
rect 9128 13379 9180 13388
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 9404 13336 9456 13388
rect 11244 13336 11296 13388
rect 11704 13336 11756 13388
rect 12624 13336 12676 13388
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 15384 13379 15436 13388
rect 15384 13345 15393 13379
rect 15393 13345 15427 13379
rect 15427 13345 15436 13379
rect 15384 13336 15436 13345
rect 16672 13336 16724 13388
rect 16948 13379 17000 13388
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 17040 13336 17092 13388
rect 26240 13404 26292 13456
rect 27252 13404 27304 13456
rect 20904 13336 20956 13388
rect 22836 13336 22888 13388
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 4160 13268 4212 13320
rect 5448 13268 5500 13320
rect 4620 13200 4672 13252
rect 3976 13132 4028 13184
rect 7196 13268 7248 13320
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 13084 13268 13136 13320
rect 13452 13268 13504 13320
rect 6000 13200 6052 13252
rect 8208 13200 8260 13252
rect 7104 13132 7156 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 9036 13200 9088 13252
rect 11520 13200 11572 13252
rect 12072 13200 12124 13252
rect 13544 13200 13596 13252
rect 16120 13268 16172 13320
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 18788 13268 18840 13320
rect 19708 13268 19760 13320
rect 9588 13132 9640 13184
rect 11244 13132 11296 13184
rect 12348 13132 12400 13184
rect 13728 13132 13780 13184
rect 15108 13132 15160 13184
rect 20168 13268 20220 13320
rect 20812 13268 20864 13320
rect 23388 13268 23440 13320
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 25872 13268 25924 13320
rect 28080 13336 28132 13388
rect 27252 13311 27304 13320
rect 27252 13277 27261 13311
rect 27261 13277 27295 13311
rect 27295 13277 27304 13311
rect 27252 13268 27304 13277
rect 34796 13268 34848 13320
rect 17960 13175 18012 13184
rect 17960 13141 17969 13175
rect 17969 13141 18003 13175
rect 18003 13141 18012 13175
rect 17960 13132 18012 13141
rect 18696 13175 18748 13184
rect 18696 13141 18705 13175
rect 18705 13141 18739 13175
rect 18739 13141 18748 13175
rect 18696 13132 18748 13141
rect 20260 13200 20312 13252
rect 20352 13200 20404 13252
rect 22744 13200 22796 13252
rect 20720 13132 20772 13184
rect 20996 13132 21048 13184
rect 23664 13132 23716 13184
rect 37280 13200 37332 13252
rect 27344 13175 27396 13184
rect 27344 13141 27353 13175
rect 27353 13141 27387 13175
rect 27387 13141 27396 13175
rect 27344 13132 27396 13141
rect 38200 13175 38252 13184
rect 38200 13141 38209 13175
rect 38209 13141 38243 13175
rect 38243 13141 38252 13175
rect 38200 13132 38252 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3332 12928 3384 12980
rect 4068 12860 4120 12912
rect 6092 12928 6144 12980
rect 6828 12860 6880 12912
rect 7932 12860 7984 12912
rect 9220 12903 9272 12912
rect 9220 12869 9229 12903
rect 9229 12869 9263 12903
rect 9263 12869 9272 12903
rect 9220 12860 9272 12869
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 2044 12588 2096 12640
rect 6000 12792 6052 12844
rect 7104 12792 7156 12844
rect 9128 12792 9180 12844
rect 14740 12928 14792 12980
rect 15108 12928 15160 12980
rect 17132 12928 17184 12980
rect 9680 12903 9732 12912
rect 9680 12869 9689 12903
rect 9689 12869 9723 12903
rect 9723 12869 9732 12903
rect 9680 12860 9732 12869
rect 10048 12860 10100 12912
rect 11244 12860 11296 12912
rect 13728 12903 13780 12912
rect 13728 12869 13737 12903
rect 13737 12869 13771 12903
rect 13771 12869 13780 12903
rect 13728 12860 13780 12869
rect 14188 12903 14240 12912
rect 14188 12869 14197 12903
rect 14197 12869 14231 12903
rect 14231 12869 14240 12903
rect 14188 12860 14240 12869
rect 18696 12903 18748 12912
rect 11704 12835 11756 12844
rect 3332 12767 3384 12776
rect 3332 12733 3341 12767
rect 3341 12733 3375 12767
rect 3375 12733 3384 12767
rect 3332 12724 3384 12733
rect 4160 12724 4212 12776
rect 5540 12724 5592 12776
rect 8668 12724 8720 12776
rect 9312 12724 9364 12776
rect 11244 12724 11296 12776
rect 8944 12656 8996 12708
rect 9956 12656 10008 12708
rect 4988 12588 5040 12640
rect 7288 12588 7340 12640
rect 7840 12588 7892 12640
rect 9128 12588 9180 12640
rect 9496 12588 9548 12640
rect 11152 12588 11204 12640
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 12624 12724 12676 12776
rect 14004 12724 14056 12776
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 14096 12656 14148 12708
rect 15016 12588 15068 12640
rect 17684 12724 17736 12776
rect 17224 12656 17276 12708
rect 18696 12869 18705 12903
rect 18705 12869 18739 12903
rect 18739 12869 18748 12903
rect 18696 12860 18748 12869
rect 19984 12928 20036 12980
rect 23940 12928 23992 12980
rect 22744 12903 22796 12912
rect 22744 12869 22753 12903
rect 22753 12869 22787 12903
rect 22787 12869 22796 12903
rect 22744 12860 22796 12869
rect 23388 12903 23440 12912
rect 23388 12869 23397 12903
rect 23397 12869 23431 12903
rect 23431 12869 23440 12903
rect 23388 12860 23440 12869
rect 18788 12724 18840 12776
rect 18972 12724 19024 12776
rect 19616 12767 19668 12776
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 21824 12792 21876 12844
rect 17316 12631 17368 12640
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 17960 12631 18012 12640
rect 17960 12597 17969 12631
rect 17969 12597 18003 12631
rect 18003 12597 18012 12631
rect 17960 12588 18012 12597
rect 20352 12656 20404 12708
rect 20444 12656 20496 12708
rect 23296 12835 23348 12844
rect 23296 12801 23305 12835
rect 23305 12801 23339 12835
rect 23339 12801 23348 12835
rect 23296 12792 23348 12801
rect 38292 12835 38344 12844
rect 38292 12801 38301 12835
rect 38301 12801 38335 12835
rect 38335 12801 38344 12835
rect 38292 12792 38344 12801
rect 19984 12588 20036 12640
rect 20628 12588 20680 12640
rect 20996 12588 21048 12640
rect 22100 12631 22152 12640
rect 22100 12597 22109 12631
rect 22109 12597 22143 12631
rect 22143 12597 22152 12631
rect 22100 12588 22152 12597
rect 22560 12588 22612 12640
rect 22836 12588 22888 12640
rect 38108 12631 38160 12640
rect 38108 12597 38117 12631
rect 38117 12597 38151 12631
rect 38151 12597 38160 12631
rect 38108 12588 38160 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3148 12384 3200 12436
rect 3332 12384 3384 12436
rect 1584 12248 1636 12300
rect 4068 12384 4120 12436
rect 4712 12384 4764 12436
rect 5448 12384 5500 12436
rect 4252 12248 4304 12300
rect 9312 12384 9364 12436
rect 10692 12384 10744 12436
rect 12716 12384 12768 12436
rect 13544 12427 13596 12436
rect 13544 12393 13553 12427
rect 13553 12393 13587 12427
rect 13587 12393 13596 12427
rect 13544 12384 13596 12393
rect 13728 12384 13780 12436
rect 16028 12359 16080 12368
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 7104 12248 7156 12300
rect 8024 12248 8076 12300
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 16028 12325 16037 12359
rect 16037 12325 16071 12359
rect 16071 12325 16080 12359
rect 16028 12316 16080 12325
rect 16580 12316 16632 12368
rect 14096 12248 14148 12300
rect 14556 12248 14608 12300
rect 16856 12248 16908 12300
rect 5356 12180 5408 12232
rect 6736 12223 6788 12232
rect 6736 12189 6745 12223
rect 6745 12189 6779 12223
rect 6779 12189 6788 12223
rect 6736 12180 6788 12189
rect 8576 12180 8628 12232
rect 4160 12112 4212 12164
rect 4252 12155 4304 12164
rect 4252 12121 4261 12155
rect 4261 12121 4295 12155
rect 4295 12121 4304 12155
rect 4252 12112 4304 12121
rect 5540 12112 5592 12164
rect 3240 12044 3292 12096
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 3516 12044 3568 12096
rect 9036 12112 9088 12164
rect 9772 12112 9824 12164
rect 10048 12112 10100 12164
rect 10232 12180 10284 12232
rect 13360 12180 13412 12232
rect 14004 12180 14056 12232
rect 11244 12112 11296 12164
rect 11428 12112 11480 12164
rect 11796 12112 11848 12164
rect 12256 12112 12308 12164
rect 12900 12112 12952 12164
rect 13912 12044 13964 12096
rect 15016 12112 15068 12164
rect 16396 12180 16448 12232
rect 18144 12384 18196 12436
rect 20536 12316 20588 12368
rect 21272 12384 21324 12436
rect 23296 12427 23348 12436
rect 23296 12393 23305 12427
rect 23305 12393 23339 12427
rect 23339 12393 23348 12427
rect 23296 12384 23348 12393
rect 20904 12248 20956 12300
rect 21916 12223 21968 12232
rect 21916 12189 21925 12223
rect 21925 12189 21959 12223
rect 21959 12189 21968 12223
rect 21916 12180 21968 12189
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 38108 12180 38160 12232
rect 16212 12112 16264 12164
rect 16672 12155 16724 12164
rect 16672 12121 16681 12155
rect 16681 12121 16715 12155
rect 16715 12121 16724 12155
rect 17224 12155 17276 12164
rect 16672 12112 16724 12121
rect 17224 12121 17233 12155
rect 17233 12121 17267 12155
rect 17267 12121 17276 12155
rect 17224 12112 17276 12121
rect 19984 12112 20036 12164
rect 20444 12155 20496 12164
rect 20444 12121 20453 12155
rect 20453 12121 20487 12155
rect 20487 12121 20496 12155
rect 20444 12112 20496 12121
rect 21272 12112 21324 12164
rect 16488 12044 16540 12096
rect 16764 12044 16816 12096
rect 20812 12044 20864 12096
rect 21088 12044 21140 12096
rect 21548 12112 21600 12164
rect 21732 12044 21784 12096
rect 22468 12044 22520 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 1952 11840 2004 11892
rect 3608 11840 3660 11892
rect 4160 11840 4212 11892
rect 1860 11815 1912 11824
rect 1860 11781 1869 11815
rect 1869 11781 1903 11815
rect 1903 11781 1912 11815
rect 1860 11772 1912 11781
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 4620 11772 4672 11824
rect 1216 11636 1268 11688
rect 1952 11636 2004 11688
rect 3516 11636 3568 11688
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 2320 11500 2372 11552
rect 3516 11500 3568 11552
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 9036 11840 9088 11892
rect 6736 11772 6788 11824
rect 7840 11772 7892 11824
rect 7012 11704 7064 11756
rect 8484 11772 8536 11824
rect 9956 11840 10008 11892
rect 10692 11772 10744 11824
rect 9864 11704 9916 11756
rect 11520 11840 11572 11892
rect 11704 11840 11756 11892
rect 14004 11840 14056 11892
rect 14648 11840 14700 11892
rect 16764 11840 16816 11892
rect 11980 11815 12032 11824
rect 11980 11781 11989 11815
rect 11989 11781 12023 11815
rect 12023 11781 12032 11815
rect 11980 11772 12032 11781
rect 12440 11772 12492 11824
rect 11428 11704 11480 11756
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 14556 11772 14608 11824
rect 14740 11772 14792 11824
rect 18604 11840 18656 11892
rect 11152 11636 11204 11688
rect 11244 11636 11296 11688
rect 17960 11772 18012 11824
rect 22100 11840 22152 11892
rect 24860 11883 24912 11892
rect 24860 11849 24869 11883
rect 24869 11849 24903 11883
rect 24903 11849 24912 11883
rect 24860 11840 24912 11849
rect 20628 11772 20680 11824
rect 20720 11772 20772 11824
rect 23112 11815 23164 11824
rect 23112 11781 23121 11815
rect 23121 11781 23155 11815
rect 23155 11781 23164 11815
rect 23112 11772 23164 11781
rect 16948 11679 17000 11688
rect 16948 11645 16957 11679
rect 16957 11645 16991 11679
rect 16991 11645 17000 11679
rect 16948 11636 17000 11645
rect 17040 11636 17092 11688
rect 20444 11679 20496 11688
rect 20444 11645 20453 11679
rect 20453 11645 20487 11679
rect 20487 11645 20496 11679
rect 21548 11704 21600 11756
rect 23572 11704 23624 11756
rect 24032 11704 24084 11756
rect 24768 11747 24820 11756
rect 24768 11713 24777 11747
rect 24777 11713 24811 11747
rect 24811 11713 24820 11747
rect 24768 11704 24820 11713
rect 38108 11704 38160 11756
rect 20444 11636 20496 11645
rect 7656 11568 7708 11620
rect 5264 11500 5316 11552
rect 5540 11500 5592 11552
rect 10416 11568 10468 11620
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 12532 11500 12584 11552
rect 13452 11500 13504 11552
rect 17132 11568 17184 11620
rect 15752 11500 15804 11552
rect 17040 11500 17092 11552
rect 17224 11500 17276 11552
rect 21180 11568 21232 11620
rect 22192 11636 22244 11688
rect 23112 11568 23164 11620
rect 21640 11500 21692 11552
rect 21732 11500 21784 11552
rect 22468 11500 22520 11552
rect 22560 11500 22612 11552
rect 26148 11500 26200 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 5724 11296 5776 11348
rect 6736 11296 6788 11348
rect 7564 11296 7616 11348
rect 7656 11296 7708 11348
rect 8024 11228 8076 11280
rect 8668 11296 8720 11348
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 10324 11296 10376 11348
rect 9220 11228 9272 11280
rect 12900 11271 12952 11280
rect 12900 11237 12909 11271
rect 12909 11237 12943 11271
rect 12943 11237 12952 11271
rect 12900 11228 12952 11237
rect 13728 11228 13780 11280
rect 3516 11160 3568 11212
rect 4252 11160 4304 11212
rect 4620 11160 4672 11212
rect 5264 11160 5316 11212
rect 5816 11160 5868 11212
rect 8392 11160 8444 11212
rect 8944 11160 8996 11212
rect 9036 11160 9088 11212
rect 8208 11092 8260 11144
rect 9680 11092 9732 11144
rect 11980 11160 12032 11212
rect 13452 11160 13504 11212
rect 14556 11160 14608 11212
rect 10600 11092 10652 11144
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 11152 11092 11204 11101
rect 12900 11092 12952 11144
rect 14004 11092 14056 11144
rect 1032 11024 1084 11076
rect 1308 11024 1360 11076
rect 4620 11067 4672 11076
rect 1768 10956 1820 11008
rect 4620 11033 4629 11067
rect 4629 11033 4663 11067
rect 4663 11033 4672 11067
rect 4620 11024 4672 11033
rect 7196 11024 7248 11076
rect 7380 11024 7432 11076
rect 11336 11024 11388 11076
rect 11888 11024 11940 11076
rect 13728 11024 13780 11076
rect 14556 11067 14608 11076
rect 12440 10956 12492 11008
rect 14556 11033 14565 11067
rect 14565 11033 14599 11067
rect 14599 11033 14608 11067
rect 14556 11024 14608 11033
rect 17960 11296 18012 11348
rect 21732 11296 21784 11348
rect 16304 11228 16356 11280
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 17040 11228 17092 11280
rect 18420 11092 18472 11144
rect 20444 11228 20496 11280
rect 24768 11296 24820 11348
rect 38108 11339 38160 11348
rect 38108 11305 38117 11339
rect 38117 11305 38151 11339
rect 38151 11305 38160 11339
rect 38108 11296 38160 11305
rect 21916 11228 21968 11280
rect 26884 11228 26936 11280
rect 22192 11160 22244 11212
rect 23296 11135 23348 11144
rect 17224 11024 17276 11076
rect 14832 10956 14884 11008
rect 19340 10956 19392 11008
rect 20628 11024 20680 11076
rect 20996 11024 21048 11076
rect 21088 11024 21140 11076
rect 23296 11101 23305 11135
rect 23305 11101 23339 11135
rect 23339 11101 23348 11135
rect 23296 11092 23348 11101
rect 26148 11135 26200 11144
rect 21916 11067 21968 11076
rect 21916 11033 21925 11067
rect 21925 11033 21959 11067
rect 21959 11033 21968 11067
rect 22836 11067 22888 11076
rect 21916 11024 21968 11033
rect 22836 11033 22845 11067
rect 22845 11033 22879 11067
rect 22879 11033 22888 11067
rect 22836 11024 22888 11033
rect 23112 11024 23164 11076
rect 26148 11101 26157 11135
rect 26157 11101 26191 11135
rect 26191 11101 26200 11135
rect 26148 11092 26200 11101
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 20536 10956 20588 11008
rect 24768 10956 24820 11008
rect 25964 10999 26016 11008
rect 25964 10965 25973 10999
rect 25973 10965 26007 10999
rect 26007 10965 26016 10999
rect 25964 10956 26016 10965
rect 26608 10999 26660 11008
rect 26608 10965 26617 10999
rect 26617 10965 26651 10999
rect 26651 10965 26660 10999
rect 26608 10956 26660 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 2320 10795 2372 10804
rect 2320 10761 2329 10795
rect 2329 10761 2363 10795
rect 2363 10761 2372 10795
rect 2320 10752 2372 10761
rect 2504 10752 2556 10804
rect 3332 10752 3384 10804
rect 6460 10752 6512 10804
rect 6644 10752 6696 10804
rect 940 10684 992 10736
rect 3424 10684 3476 10736
rect 6828 10684 6880 10736
rect 3056 10616 3108 10668
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 7748 10684 7800 10736
rect 7288 10616 7340 10668
rect 8024 10684 8076 10736
rect 8392 10684 8444 10736
rect 10600 10684 10652 10736
rect 11888 10752 11940 10804
rect 12164 10752 12216 10804
rect 12256 10684 12308 10736
rect 13268 10684 13320 10736
rect 15660 10684 15712 10736
rect 10140 10616 10192 10668
rect 10232 10616 10284 10668
rect 11336 10616 11388 10668
rect 11060 10548 11112 10600
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 12072 10548 12124 10600
rect 12348 10548 12400 10600
rect 3792 10480 3844 10532
rect 5264 10412 5316 10464
rect 7840 10480 7892 10532
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 7104 10412 7156 10464
rect 7288 10412 7340 10464
rect 7472 10412 7524 10464
rect 9680 10412 9732 10464
rect 10508 10412 10560 10464
rect 10784 10412 10836 10464
rect 13728 10412 13780 10464
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 14280 10548 14332 10600
rect 14832 10548 14884 10600
rect 14832 10412 14884 10464
rect 18880 10752 18932 10804
rect 24124 10795 24176 10804
rect 24124 10761 24133 10795
rect 24133 10761 24167 10795
rect 24167 10761 24176 10795
rect 24124 10752 24176 10761
rect 16764 10616 16816 10668
rect 17500 10684 17552 10736
rect 18512 10727 18564 10736
rect 18512 10693 18521 10727
rect 18521 10693 18555 10727
rect 18555 10693 18564 10727
rect 18512 10684 18564 10693
rect 19432 10727 19484 10736
rect 19432 10693 19441 10727
rect 19441 10693 19475 10727
rect 19475 10693 19484 10727
rect 19432 10684 19484 10693
rect 20812 10684 20864 10736
rect 21180 10727 21232 10736
rect 21180 10693 21189 10727
rect 21189 10693 21223 10727
rect 21223 10693 21232 10727
rect 21180 10684 21232 10693
rect 21272 10684 21324 10736
rect 22008 10684 22060 10736
rect 17316 10616 17368 10668
rect 21548 10616 21600 10668
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 16948 10548 17000 10600
rect 18512 10548 18564 10600
rect 18880 10548 18932 10600
rect 19064 10548 19116 10600
rect 19984 10548 20036 10600
rect 21088 10548 21140 10600
rect 22100 10548 22152 10600
rect 25872 10684 25924 10736
rect 25964 10659 26016 10668
rect 25964 10625 25973 10659
rect 25973 10625 26007 10659
rect 26007 10625 26016 10659
rect 25964 10616 26016 10625
rect 24216 10548 24268 10600
rect 26608 10548 26660 10600
rect 33048 10616 33100 10668
rect 38108 10548 38160 10600
rect 16488 10480 16540 10532
rect 23112 10480 23164 10532
rect 17500 10412 17552 10464
rect 20996 10412 21048 10464
rect 21180 10412 21232 10464
rect 22928 10412 22980 10464
rect 24492 10412 24544 10464
rect 30932 10455 30984 10464
rect 30932 10421 30941 10455
rect 30941 10421 30975 10455
rect 30975 10421 30984 10455
rect 30932 10412 30984 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2964 10208 3016 10260
rect 5632 10208 5684 10260
rect 6644 10208 6696 10260
rect 16396 10208 16448 10260
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 18236 10208 18288 10260
rect 19708 10208 19760 10260
rect 22284 10208 22336 10260
rect 22928 10208 22980 10260
rect 8392 10140 8444 10192
rect 11336 10140 11388 10192
rect 11888 10140 11940 10192
rect 13452 10140 13504 10192
rect 15844 10140 15896 10192
rect 16856 10140 16908 10192
rect 19064 10140 19116 10192
rect 2596 10072 2648 10124
rect 5908 10072 5960 10124
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 7472 10072 7524 10124
rect 7656 10072 7708 10124
rect 7748 10072 7800 10124
rect 11060 10072 11112 10124
rect 14924 10072 14976 10124
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 17408 10072 17460 10124
rect 18696 10115 18748 10124
rect 18696 10081 18705 10115
rect 18705 10081 18739 10115
rect 18739 10081 18748 10115
rect 19432 10140 19484 10192
rect 20260 10140 20312 10192
rect 18696 10072 18748 10081
rect 19892 10072 19944 10124
rect 19984 10072 20036 10124
rect 21640 10072 21692 10124
rect 24216 10072 24268 10124
rect 6644 10004 6696 10056
rect 1952 9979 2004 9988
rect 1952 9945 1961 9979
rect 1961 9945 1995 9979
rect 1995 9945 2004 9979
rect 1952 9936 2004 9945
rect 3516 9936 3568 9988
rect 5908 9936 5960 9988
rect 5080 9868 5132 9920
rect 5264 9868 5316 9920
rect 6092 9868 6144 9920
rect 11152 9936 11204 9988
rect 16212 10004 16264 10056
rect 16672 10004 16724 10056
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 19156 10004 19208 10056
rect 24768 10047 24820 10056
rect 24768 10013 24777 10047
rect 24777 10013 24811 10047
rect 24811 10013 24820 10047
rect 24768 10004 24820 10013
rect 26056 10047 26108 10056
rect 26056 10013 26065 10047
rect 26065 10013 26099 10047
rect 26099 10013 26108 10047
rect 26056 10004 26108 10013
rect 34520 10072 34572 10124
rect 37188 10004 37240 10056
rect 12164 9979 12216 9988
rect 12164 9945 12173 9979
rect 12173 9945 12207 9979
rect 12207 9945 12216 9979
rect 12164 9936 12216 9945
rect 12808 9936 12860 9988
rect 13728 9936 13780 9988
rect 16396 9936 16448 9988
rect 18604 9936 18656 9988
rect 8484 9868 8536 9920
rect 9680 9868 9732 9920
rect 9772 9868 9824 9920
rect 10508 9868 10560 9920
rect 13084 9868 13136 9920
rect 15936 9868 15988 9920
rect 19524 9936 19576 9988
rect 19892 9936 19944 9988
rect 21824 9979 21876 9988
rect 20536 9868 20588 9920
rect 21824 9945 21833 9979
rect 21833 9945 21867 9979
rect 21867 9945 21876 9979
rect 21824 9936 21876 9945
rect 22100 9936 22152 9988
rect 23848 9979 23900 9988
rect 22744 9868 22796 9920
rect 23848 9945 23857 9979
rect 23857 9945 23891 9979
rect 23891 9945 23900 9979
rect 23848 9936 23900 9945
rect 28264 9936 28316 9988
rect 33140 9936 33192 9988
rect 34428 9936 34480 9988
rect 25964 9868 26016 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 5908 9664 5960 9716
rect 10508 9664 10560 9716
rect 15200 9664 15252 9716
rect 17408 9664 17460 9716
rect 3516 9596 3568 9648
rect 8024 9596 8076 9648
rect 9588 9596 9640 9648
rect 13452 9596 13504 9648
rect 14188 9596 14240 9648
rect 5908 9528 5960 9580
rect 6552 9528 6604 9580
rect 2504 9460 2556 9512
rect 2228 9324 2280 9376
rect 2596 9324 2648 9376
rect 3424 9324 3476 9376
rect 3884 9324 3936 9376
rect 5540 9460 5592 9512
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 6552 9435 6604 9444
rect 6552 9401 6561 9435
rect 6561 9401 6595 9435
rect 6595 9401 6604 9435
rect 6552 9392 6604 9401
rect 4712 9324 4764 9376
rect 5172 9324 5224 9376
rect 6920 9460 6972 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7840 9460 7892 9512
rect 8116 9460 8168 9512
rect 9772 9528 9824 9580
rect 10508 9528 10560 9580
rect 11152 9528 11204 9580
rect 16028 9596 16080 9648
rect 17960 9664 18012 9716
rect 17776 9596 17828 9648
rect 20352 9664 20404 9716
rect 21088 9664 21140 9716
rect 30932 9664 30984 9716
rect 7840 9324 7892 9376
rect 11796 9460 11848 9512
rect 12164 9503 12216 9512
rect 10416 9392 10468 9444
rect 11704 9392 11756 9444
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 10140 9324 10192 9376
rect 11796 9324 11848 9376
rect 13176 9392 13228 9444
rect 14004 9460 14056 9512
rect 14280 9460 14332 9512
rect 15384 9460 15436 9512
rect 16488 9528 16540 9580
rect 21272 9596 21324 9648
rect 22376 9596 22428 9648
rect 22744 9639 22796 9648
rect 22744 9605 22753 9639
rect 22753 9605 22787 9639
rect 22787 9605 22796 9639
rect 22744 9596 22796 9605
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 16396 9392 16448 9444
rect 16856 9392 16908 9444
rect 17408 9460 17460 9512
rect 19156 9528 19208 9580
rect 21824 9528 21876 9580
rect 21916 9528 21968 9580
rect 23112 9528 23164 9580
rect 24032 9528 24084 9580
rect 24492 9571 24544 9580
rect 24492 9537 24501 9571
rect 24501 9537 24535 9571
rect 24535 9537 24544 9571
rect 24492 9528 24544 9537
rect 24584 9528 24636 9580
rect 18052 9460 18104 9512
rect 19892 9503 19944 9512
rect 17776 9392 17828 9444
rect 19892 9469 19901 9503
rect 19901 9469 19935 9503
rect 19935 9469 19944 9503
rect 19892 9460 19944 9469
rect 20536 9460 20588 9512
rect 18880 9392 18932 9444
rect 23204 9392 23256 9444
rect 14464 9324 14516 9376
rect 15752 9324 15804 9376
rect 15936 9324 15988 9376
rect 19892 9324 19944 9376
rect 22100 9367 22152 9376
rect 22100 9333 22109 9367
rect 22109 9333 22143 9367
rect 22143 9333 22152 9367
rect 22100 9324 22152 9333
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2596 9163 2648 9172
rect 2596 9129 2605 9163
rect 2605 9129 2639 9163
rect 2639 9129 2648 9163
rect 2596 9120 2648 9129
rect 2688 9120 2740 9172
rect 2136 9052 2188 9104
rect 3608 9052 3660 9104
rect 4620 9052 4672 9104
rect 7748 9120 7800 9172
rect 11520 9120 11572 9172
rect 5908 9052 5960 9104
rect 7564 9052 7616 9104
rect 4712 9027 4764 9036
rect 1492 8916 1544 8968
rect 2504 8916 2556 8968
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 2780 8916 2832 8925
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 6460 9027 6512 9036
rect 6460 8993 6469 9027
rect 6469 8993 6503 9027
rect 6503 8993 6512 9027
rect 6460 8984 6512 8993
rect 6552 8984 6604 9036
rect 4896 8916 4948 8968
rect 4620 8848 4672 8900
rect 5908 8916 5960 8968
rect 8024 8916 8076 8968
rect 9864 8916 9916 8968
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 5632 8848 5684 8900
rect 6736 8848 6788 8900
rect 7748 8848 7800 8900
rect 10416 8984 10468 9036
rect 10968 8984 11020 9036
rect 11612 8984 11664 9036
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 14924 8984 14976 9036
rect 16488 9052 16540 9104
rect 18512 9052 18564 9104
rect 18696 9120 18748 9172
rect 18972 9120 19024 9172
rect 19984 9120 20036 9172
rect 20720 9163 20772 9172
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 23848 9163 23900 9172
rect 23848 9129 23857 9163
rect 23857 9129 23891 9163
rect 23891 9129 23900 9163
rect 23848 9120 23900 9129
rect 24584 9163 24636 9172
rect 24584 9129 24593 9163
rect 24593 9129 24627 9163
rect 24627 9129 24636 9163
rect 24584 9120 24636 9129
rect 25504 9120 25556 9172
rect 18880 9052 18932 9104
rect 18788 8984 18840 9036
rect 22652 9052 22704 9104
rect 19984 9027 20036 9036
rect 19984 8993 19993 9027
rect 19993 8993 20027 9027
rect 20027 8993 20036 9027
rect 19984 8984 20036 8993
rect 20904 8984 20956 9036
rect 23388 8984 23440 9036
rect 12348 8916 12400 8968
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 13728 8916 13780 8968
rect 14004 8916 14056 8968
rect 16212 8916 16264 8968
rect 17776 8916 17828 8968
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 20352 8916 20404 8968
rect 8760 8780 8812 8832
rect 9956 8823 10008 8832
rect 9956 8789 9965 8823
rect 9965 8789 9999 8823
rect 9999 8789 10008 8823
rect 9956 8780 10008 8789
rect 14556 8891 14608 8900
rect 14556 8857 14565 8891
rect 14565 8857 14599 8891
rect 14599 8857 14608 8891
rect 14556 8848 14608 8857
rect 15200 8848 15252 8900
rect 12532 8780 12584 8832
rect 16580 8848 16632 8900
rect 18052 8891 18104 8900
rect 15936 8780 15988 8832
rect 18052 8857 18061 8891
rect 18061 8857 18095 8891
rect 18095 8857 18104 8891
rect 18052 8848 18104 8857
rect 18144 8891 18196 8900
rect 18144 8857 18153 8891
rect 18153 8857 18187 8891
rect 18187 8857 18196 8891
rect 18144 8848 18196 8857
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 17592 8780 17644 8832
rect 18880 8780 18932 8832
rect 19340 8780 19392 8832
rect 20812 8848 20864 8900
rect 21180 8848 21232 8900
rect 21456 8891 21508 8900
rect 21456 8857 21465 8891
rect 21465 8857 21499 8891
rect 21499 8857 21508 8891
rect 21456 8848 21508 8857
rect 21732 8848 21784 8900
rect 21916 8780 21968 8832
rect 22744 8916 22796 8968
rect 23940 8916 23992 8968
rect 25228 8959 25280 8968
rect 25228 8925 25237 8959
rect 25237 8925 25271 8959
rect 25271 8925 25280 8959
rect 25228 8916 25280 8925
rect 30748 8916 30800 8968
rect 22560 8780 22612 8832
rect 25320 8823 25372 8832
rect 25320 8789 25329 8823
rect 25329 8789 25363 8823
rect 25363 8789 25372 8823
rect 25320 8780 25372 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1400 8576 1452 8628
rect 2872 8576 2924 8628
rect 7748 8576 7800 8628
rect 2964 8508 3016 8560
rect 4712 8508 4764 8560
rect 5540 8508 5592 8560
rect 3976 8440 4028 8492
rect 9404 8576 9456 8628
rect 9956 8576 10008 8628
rect 13268 8576 13320 8628
rect 13912 8576 13964 8628
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 17868 8576 17920 8628
rect 19708 8576 19760 8628
rect 8484 8508 8536 8560
rect 9220 8508 9272 8560
rect 2228 8372 2280 8424
rect 1308 8304 1360 8356
rect 4988 8372 5040 8424
rect 5540 8372 5592 8424
rect 5724 8372 5776 8424
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 9312 8372 9364 8424
rect 10416 8440 10468 8492
rect 12348 8508 12400 8560
rect 12992 8508 13044 8560
rect 13544 8508 13596 8560
rect 14740 8551 14792 8560
rect 14740 8517 14749 8551
rect 14749 8517 14783 8551
rect 14783 8517 14792 8551
rect 14740 8508 14792 8517
rect 15108 8508 15160 8560
rect 10784 8440 10836 8492
rect 11152 8440 11204 8492
rect 11704 8440 11756 8492
rect 10876 8372 10928 8424
rect 11244 8372 11296 8424
rect 12716 8372 12768 8424
rect 14464 8440 14516 8492
rect 18052 8508 18104 8560
rect 18604 8508 18656 8560
rect 16764 8440 16816 8492
rect 14096 8372 14148 8424
rect 15108 8372 15160 8424
rect 15568 8372 15620 8424
rect 15752 8372 15804 8424
rect 3700 8304 3752 8356
rect 7380 8304 7432 8356
rect 5724 8236 5776 8288
rect 6552 8236 6604 8288
rect 9128 8304 9180 8356
rect 10508 8304 10560 8356
rect 13728 8304 13780 8356
rect 17592 8440 17644 8492
rect 20996 8576 21048 8628
rect 22100 8576 22152 8628
rect 21364 8551 21416 8560
rect 21364 8517 21373 8551
rect 21373 8517 21407 8551
rect 21407 8517 21416 8551
rect 21364 8508 21416 8517
rect 21456 8508 21508 8560
rect 33048 8576 33100 8628
rect 20720 8440 20772 8492
rect 21088 8440 21140 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 18236 8372 18288 8424
rect 18512 8372 18564 8424
rect 18604 8415 18656 8424
rect 18604 8381 18613 8415
rect 18613 8381 18647 8415
rect 18647 8381 18656 8415
rect 18604 8372 18656 8381
rect 19064 8372 19116 8424
rect 19800 8372 19852 8424
rect 20352 8372 20404 8424
rect 20904 8372 20956 8424
rect 20996 8372 21048 8424
rect 23388 8440 23440 8492
rect 25044 8483 25096 8492
rect 25044 8449 25053 8483
rect 25053 8449 25087 8483
rect 25087 8449 25096 8483
rect 25044 8440 25096 8449
rect 38292 8483 38344 8492
rect 20536 8304 20588 8356
rect 22376 8304 22428 8356
rect 24860 8304 24912 8356
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 26148 8304 26200 8356
rect 34428 8304 34480 8356
rect 9312 8236 9364 8288
rect 10232 8236 10284 8288
rect 10416 8236 10468 8288
rect 11244 8236 11296 8288
rect 15200 8236 15252 8288
rect 16488 8236 16540 8288
rect 24768 8236 24820 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1676 8032 1728 8084
rect 4528 7964 4580 8016
rect 5632 7964 5684 8016
rect 940 7896 992 7948
rect 3792 7896 3844 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4988 7896 5040 7948
rect 13544 8032 13596 8084
rect 14188 8032 14240 8084
rect 16396 8032 16448 8084
rect 18052 8032 18104 8084
rect 18236 8032 18288 8084
rect 7656 8007 7708 8016
rect 7656 7973 7665 8007
rect 7665 7973 7699 8007
rect 7699 7973 7708 8007
rect 7656 7964 7708 7973
rect 6644 7896 6696 7948
rect 8300 7896 8352 7948
rect 8852 7896 8904 7948
rect 9128 7939 9180 7948
rect 9128 7905 9137 7939
rect 9137 7905 9171 7939
rect 9171 7905 9180 7939
rect 9128 7896 9180 7905
rect 10968 7964 11020 8016
rect 16028 8007 16080 8016
rect 16028 7973 16037 8007
rect 16037 7973 16071 8007
rect 16071 7973 16080 8007
rect 16028 7964 16080 7973
rect 11152 7896 11204 7948
rect 11704 7896 11756 7948
rect 13636 7896 13688 7948
rect 15200 7939 15252 7948
rect 15200 7905 15209 7939
rect 15209 7905 15243 7939
rect 15243 7905 15252 7939
rect 15200 7896 15252 7905
rect 17500 7896 17552 7948
rect 17592 7939 17644 7948
rect 17592 7905 17601 7939
rect 17601 7905 17635 7939
rect 17635 7905 17644 7939
rect 17592 7896 17644 7905
rect 17776 7896 17828 7948
rect 18420 7964 18472 8016
rect 20076 7964 20128 8016
rect 20260 8032 20312 8084
rect 20720 8032 20772 8084
rect 20812 8032 20864 8084
rect 31392 8075 31444 8084
rect 31392 8041 31401 8075
rect 31401 8041 31435 8075
rect 31435 8041 31444 8075
rect 31392 8032 31444 8041
rect 5724 7828 5776 7880
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6460 7760 6512 7812
rect 4988 7692 5040 7744
rect 8208 7760 8260 7812
rect 11060 7828 11112 7880
rect 16488 7828 16540 7880
rect 19800 7896 19852 7948
rect 20352 7939 20404 7948
rect 20352 7905 20361 7939
rect 20361 7905 20395 7939
rect 20395 7905 20404 7939
rect 20352 7896 20404 7905
rect 20720 7896 20772 7948
rect 20812 7939 20864 7948
rect 20812 7905 20821 7939
rect 20821 7905 20855 7939
rect 20855 7905 20864 7939
rect 20812 7896 20864 7905
rect 21180 7896 21232 7948
rect 21824 7896 21876 7948
rect 24032 7896 24084 7948
rect 18328 7828 18380 7880
rect 20076 7828 20128 7880
rect 20168 7828 20220 7880
rect 22652 7871 22704 7880
rect 22652 7837 22661 7871
rect 22661 7837 22695 7871
rect 22695 7837 22704 7871
rect 22652 7828 22704 7837
rect 23204 7828 23256 7880
rect 23388 7828 23440 7880
rect 34428 7828 34480 7880
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 9312 7760 9364 7812
rect 9404 7803 9456 7812
rect 9404 7769 9413 7803
rect 9413 7769 9447 7803
rect 9447 7769 9456 7803
rect 9404 7760 9456 7769
rect 10968 7760 11020 7812
rect 8392 7692 8444 7744
rect 8668 7692 8720 7744
rect 14556 7692 14608 7744
rect 16580 7692 16632 7744
rect 17868 7760 17920 7812
rect 20352 7760 20404 7812
rect 17500 7692 17552 7744
rect 17960 7692 18012 7744
rect 20168 7692 20220 7744
rect 21640 7803 21692 7812
rect 21640 7769 21649 7803
rect 21649 7769 21683 7803
rect 21683 7769 21692 7803
rect 21640 7760 21692 7769
rect 21824 7760 21876 7812
rect 22560 7692 22612 7744
rect 38016 7692 38068 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4804 7488 4856 7540
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 5356 7488 5408 7540
rect 5816 7488 5868 7540
rect 8392 7488 8444 7540
rect 9404 7488 9456 7540
rect 13176 7488 13228 7540
rect 14096 7488 14148 7540
rect 18328 7488 18380 7540
rect 5908 7420 5960 7472
rect 8576 7463 8628 7472
rect 8576 7429 8585 7463
rect 8585 7429 8619 7463
rect 8619 7429 8628 7463
rect 8576 7420 8628 7429
rect 12072 7420 12124 7472
rect 12624 7420 12676 7472
rect 13820 7420 13872 7472
rect 15384 7420 15436 7472
rect 18420 7420 18472 7472
rect 20904 7488 20956 7540
rect 21640 7488 21692 7540
rect 23020 7488 23072 7540
rect 25228 7531 25280 7540
rect 25228 7497 25237 7531
rect 25237 7497 25271 7531
rect 25271 7497 25280 7531
rect 25228 7488 25280 7497
rect 19708 7420 19760 7472
rect 20444 7420 20496 7472
rect 20628 7463 20680 7472
rect 20628 7429 20637 7463
rect 20637 7429 20671 7463
rect 20671 7429 20680 7463
rect 20628 7420 20680 7429
rect 20996 7420 21048 7472
rect 21272 7420 21324 7472
rect 1400 7352 1452 7404
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5264 7352 5316 7404
rect 5540 7352 5592 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 6644 7352 6696 7404
rect 8116 7352 8168 7404
rect 4068 7284 4120 7336
rect 5080 7284 5132 7336
rect 6920 7284 6972 7336
rect 10048 7352 10100 7404
rect 10416 7352 10468 7404
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 14188 7395 14240 7404
rect 10692 7352 10744 7361
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 8576 7284 8628 7336
rect 11244 7284 11296 7336
rect 11612 7284 11664 7336
rect 14924 7284 14976 7336
rect 15292 7284 15344 7336
rect 17316 7327 17368 7336
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 17776 7327 17828 7336
rect 17776 7293 17785 7327
rect 17785 7293 17819 7327
rect 17819 7293 17828 7327
rect 17776 7284 17828 7293
rect 18328 7284 18380 7336
rect 19156 7284 19208 7336
rect 19708 7284 19760 7336
rect 19800 7284 19852 7336
rect 20260 7284 20312 7336
rect 21272 7284 21324 7336
rect 24216 7352 24268 7404
rect 25044 7352 25096 7404
rect 23388 7284 23440 7336
rect 24860 7327 24912 7336
rect 24860 7293 24869 7327
rect 24869 7293 24903 7327
rect 24903 7293 24912 7327
rect 24860 7284 24912 7293
rect 4804 7148 4856 7200
rect 4988 7148 5040 7200
rect 8300 7148 8352 7200
rect 19064 7216 19116 7268
rect 9864 7148 9916 7200
rect 12900 7148 12952 7200
rect 16396 7148 16448 7200
rect 16488 7148 16540 7200
rect 18512 7148 18564 7200
rect 18696 7148 18748 7200
rect 21824 7216 21876 7268
rect 23480 7148 23532 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2044 6944 2096 6996
rect 6000 6944 6052 6996
rect 7196 6944 7248 6996
rect 7564 6944 7616 6996
rect 7656 6987 7708 6996
rect 7656 6953 7665 6987
rect 7665 6953 7699 6987
rect 7699 6953 7708 6987
rect 7656 6944 7708 6953
rect 8208 6944 8260 6996
rect 23204 6944 23256 6996
rect 3332 6851 3384 6860
rect 3332 6817 3341 6851
rect 3341 6817 3375 6851
rect 3375 6817 3384 6851
rect 3332 6808 3384 6817
rect 3884 6808 3936 6860
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 4620 6808 4672 6860
rect 6552 6808 6604 6860
rect 5908 6783 5960 6792
rect 5908 6749 5917 6783
rect 5917 6749 5951 6783
rect 5951 6749 5960 6783
rect 5908 6740 5960 6749
rect 8208 6740 8260 6792
rect 8760 6876 8812 6928
rect 9680 6876 9732 6928
rect 8852 6808 8904 6860
rect 9772 6808 9824 6860
rect 9036 6740 9088 6792
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 9680 6740 9732 6792
rect 21640 6876 21692 6928
rect 14004 6808 14056 6860
rect 14188 6808 14240 6860
rect 14740 6808 14792 6860
rect 15292 6808 15344 6860
rect 16488 6808 16540 6860
rect 17132 6808 17184 6860
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 4620 6672 4672 6724
rect 4988 6715 5040 6724
rect 4988 6681 4997 6715
rect 4997 6681 5031 6715
rect 5031 6681 5040 6715
rect 4988 6672 5040 6681
rect 8116 6672 8168 6724
rect 10324 6715 10376 6724
rect 10324 6681 10333 6715
rect 10333 6681 10367 6715
rect 10367 6681 10376 6715
rect 10324 6672 10376 6681
rect 12716 6672 12768 6724
rect 12900 6672 12952 6724
rect 13820 6672 13872 6724
rect 15108 6715 15160 6724
rect 15108 6681 15117 6715
rect 15117 6681 15151 6715
rect 15151 6681 15160 6715
rect 15108 6672 15160 6681
rect 17132 6672 17184 6724
rect 17316 6672 17368 6724
rect 17592 6672 17644 6724
rect 7564 6604 7616 6656
rect 9588 6604 9640 6656
rect 11060 6604 11112 6656
rect 11336 6604 11388 6656
rect 11888 6604 11940 6656
rect 13360 6604 13412 6656
rect 15200 6604 15252 6656
rect 19156 6808 19208 6860
rect 19892 6808 19944 6860
rect 19340 6740 19392 6792
rect 20260 6740 20312 6792
rect 23388 6851 23440 6860
rect 18236 6715 18288 6724
rect 18236 6681 18245 6715
rect 18245 6681 18279 6715
rect 18279 6681 18288 6715
rect 18236 6672 18288 6681
rect 18512 6672 18564 6724
rect 18880 6672 18932 6724
rect 19340 6604 19392 6656
rect 19708 6672 19760 6724
rect 22652 6740 22704 6792
rect 23388 6817 23397 6851
rect 23397 6817 23431 6851
rect 23431 6817 23440 6851
rect 23388 6808 23440 6817
rect 23480 6740 23532 6792
rect 23572 6783 23624 6792
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 24676 6740 24728 6792
rect 21364 6672 21416 6724
rect 21180 6604 21232 6656
rect 21824 6647 21876 6656
rect 21824 6613 21833 6647
rect 21833 6613 21867 6647
rect 21867 6613 21876 6647
rect 21824 6604 21876 6613
rect 22008 6604 22060 6656
rect 22192 6604 22244 6656
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 5908 6400 5960 6452
rect 6368 6332 6420 6384
rect 2320 6060 2372 6112
rect 2412 6060 2464 6112
rect 11888 6400 11940 6452
rect 7196 6375 7248 6384
rect 7196 6341 7205 6375
rect 7205 6341 7239 6375
rect 7239 6341 7248 6375
rect 7196 6332 7248 6341
rect 9036 6332 9088 6384
rect 6828 6264 6880 6316
rect 9312 6332 9364 6384
rect 9404 6375 9456 6384
rect 9404 6341 9413 6375
rect 9413 6341 9447 6375
rect 9447 6341 9456 6375
rect 9404 6332 9456 6341
rect 9864 6332 9916 6384
rect 11428 6332 11480 6384
rect 17592 6400 17644 6452
rect 13084 6264 13136 6316
rect 6552 6128 6604 6180
rect 8208 6196 8260 6248
rect 9956 6196 10008 6248
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 11244 6196 11296 6248
rect 11612 6196 11664 6248
rect 12348 6196 12400 6248
rect 14924 6332 14976 6384
rect 17224 6332 17276 6384
rect 20628 6400 20680 6452
rect 20720 6400 20772 6452
rect 21180 6400 21232 6452
rect 22468 6400 22520 6452
rect 22560 6400 22612 6452
rect 23572 6400 23624 6452
rect 30380 6400 30432 6452
rect 38108 6443 38160 6452
rect 38108 6409 38117 6443
rect 38117 6409 38151 6443
rect 38151 6409 38160 6443
rect 38108 6400 38160 6409
rect 18604 6332 18656 6384
rect 18788 6375 18840 6384
rect 18788 6341 18797 6375
rect 18797 6341 18831 6375
rect 18831 6341 18840 6375
rect 18788 6332 18840 6341
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 17316 6264 17368 6316
rect 18236 6307 18288 6316
rect 18236 6273 18245 6307
rect 18245 6273 18279 6307
rect 18279 6273 18288 6307
rect 18236 6264 18288 6273
rect 18512 6264 18564 6316
rect 19800 6332 19852 6384
rect 20536 6332 20588 6384
rect 21456 6332 21508 6384
rect 21088 6264 21140 6316
rect 21916 6332 21968 6384
rect 21732 6264 21784 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 15200 6196 15252 6248
rect 16488 6196 16540 6248
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 18328 6196 18380 6248
rect 18972 6196 19024 6248
rect 20628 6196 20680 6248
rect 24400 6332 24452 6384
rect 22928 6264 22980 6316
rect 23296 6307 23348 6316
rect 23296 6273 23305 6307
rect 23305 6273 23339 6307
rect 23339 6273 23348 6307
rect 23296 6264 23348 6273
rect 23940 6307 23992 6316
rect 23940 6273 23949 6307
rect 23949 6273 23983 6307
rect 23983 6273 23992 6307
rect 23940 6264 23992 6273
rect 26148 6307 26200 6316
rect 22836 6196 22888 6248
rect 26148 6273 26157 6307
rect 26157 6273 26191 6307
rect 26191 6273 26200 6307
rect 26148 6264 26200 6273
rect 26424 6264 26476 6316
rect 34060 6264 34112 6316
rect 38292 6307 38344 6316
rect 38292 6273 38301 6307
rect 38301 6273 38335 6307
rect 38335 6273 38344 6307
rect 38292 6264 38344 6273
rect 28448 6196 28500 6248
rect 4896 6060 4948 6112
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 10876 6060 10928 6112
rect 11060 6060 11112 6112
rect 13360 6060 13412 6112
rect 16580 6060 16632 6112
rect 17224 6060 17276 6112
rect 18604 6060 18656 6112
rect 19156 6060 19208 6112
rect 20352 6060 20404 6112
rect 21824 6128 21876 6180
rect 22008 6060 22060 6112
rect 25596 6060 25648 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3424 5856 3476 5908
rect 1584 5720 1636 5772
rect 2044 5720 2096 5772
rect 4988 5720 5040 5772
rect 6460 5856 6512 5908
rect 5632 5788 5684 5840
rect 8392 5856 8444 5908
rect 11888 5856 11940 5908
rect 13084 5856 13136 5908
rect 20720 5856 20772 5908
rect 21640 5856 21692 5908
rect 24860 5899 24912 5908
rect 24860 5865 24869 5899
rect 24869 5865 24903 5899
rect 24903 5865 24912 5899
rect 24860 5856 24912 5865
rect 26424 5899 26476 5908
rect 26424 5865 26433 5899
rect 26433 5865 26467 5899
rect 26467 5865 26476 5899
rect 26424 5856 26476 5865
rect 8116 5788 8168 5840
rect 10416 5788 10468 5840
rect 10600 5831 10652 5840
rect 10600 5797 10609 5831
rect 10609 5797 10643 5831
rect 10643 5797 10652 5831
rect 10600 5788 10652 5797
rect 10876 5788 10928 5840
rect 7196 5720 7248 5772
rect 11244 5763 11296 5772
rect 11244 5729 11253 5763
rect 11253 5729 11287 5763
rect 11287 5729 11296 5763
rect 11244 5720 11296 5729
rect 11612 5720 11664 5772
rect 13268 5788 13320 5840
rect 17132 5788 17184 5840
rect 18604 5788 18656 5840
rect 19432 5788 19484 5840
rect 20260 5788 20312 5840
rect 14648 5720 14700 5772
rect 17960 5720 18012 5772
rect 5540 5652 5592 5704
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 8576 5652 8628 5704
rect 10140 5652 10192 5704
rect 10600 5652 10652 5704
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 16764 5652 16816 5704
rect 18512 5720 18564 5772
rect 20904 5720 20956 5772
rect 18328 5652 18380 5704
rect 18696 5652 18748 5704
rect 19524 5652 19576 5704
rect 3332 5516 3384 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 4528 5584 4580 5636
rect 7196 5584 7248 5636
rect 7564 5584 7616 5636
rect 9772 5584 9824 5636
rect 3424 5516 3476 5525
rect 8116 5516 8168 5568
rect 8392 5516 8444 5568
rect 11888 5516 11940 5568
rect 14464 5584 14516 5636
rect 15016 5584 15068 5636
rect 15936 5584 15988 5636
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 18512 5584 18564 5636
rect 20352 5652 20404 5704
rect 21088 5652 21140 5704
rect 21548 5652 21600 5704
rect 21732 5652 21784 5704
rect 23664 5788 23716 5840
rect 25044 5788 25096 5840
rect 22468 5695 22520 5704
rect 22468 5661 22477 5695
rect 22477 5661 22511 5695
rect 22511 5661 22520 5695
rect 22468 5652 22520 5661
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 16028 5559 16080 5568
rect 16028 5525 16037 5559
rect 16037 5525 16071 5559
rect 16071 5525 16080 5559
rect 16028 5516 16080 5525
rect 16120 5516 16172 5568
rect 16764 5516 16816 5568
rect 21456 5516 21508 5568
rect 21824 5516 21876 5568
rect 22376 5516 22428 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3884 5244 3936 5296
rect 6828 5312 6880 5364
rect 4436 5244 4488 5296
rect 4620 5244 4672 5296
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 9772 5312 9824 5364
rect 8576 5176 8628 5228
rect 9956 5244 10008 5296
rect 14648 5287 14700 5296
rect 14648 5253 14657 5287
rect 14657 5253 14691 5287
rect 14691 5253 14700 5287
rect 14648 5244 14700 5253
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 2688 5108 2740 5160
rect 5172 5108 5224 5160
rect 6276 5108 6328 5160
rect 6644 5108 6696 5160
rect 7840 5108 7892 5160
rect 5724 5040 5776 5092
rect 10784 5176 10836 5228
rect 11244 5176 11296 5228
rect 17592 5312 17644 5364
rect 16764 5176 16816 5228
rect 11704 5151 11756 5160
rect 4528 4972 4580 5024
rect 5264 4972 5316 5024
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 11152 5083 11204 5092
rect 11152 5049 11161 5083
rect 11161 5049 11195 5083
rect 11195 5049 11204 5083
rect 11152 5040 11204 5049
rect 8944 4972 8996 4981
rect 9680 4972 9732 5024
rect 11704 5117 11713 5151
rect 11713 5117 11747 5151
rect 11747 5117 11756 5151
rect 11704 5108 11756 5117
rect 15844 5108 15896 5160
rect 15936 5040 15988 5092
rect 16580 5040 16632 5092
rect 20628 5312 20680 5364
rect 18512 5287 18564 5296
rect 18512 5253 18521 5287
rect 18521 5253 18555 5287
rect 18555 5253 18564 5287
rect 18512 5244 18564 5253
rect 18696 5244 18748 5296
rect 19064 5287 19116 5296
rect 19064 5253 19073 5287
rect 19073 5253 19107 5287
rect 19107 5253 19116 5287
rect 19064 5244 19116 5253
rect 19156 5244 19208 5296
rect 19708 5244 19760 5296
rect 20444 5176 20496 5228
rect 17224 5151 17276 5160
rect 17224 5117 17233 5151
rect 17233 5117 17267 5151
rect 17267 5117 17276 5151
rect 17224 5108 17276 5117
rect 12164 4972 12216 5024
rect 13360 4972 13412 5024
rect 15292 4972 15344 5024
rect 16856 4972 16908 5024
rect 17776 5083 17828 5092
rect 17776 5049 17785 5083
rect 17785 5049 17819 5083
rect 17819 5049 17828 5083
rect 19432 5108 19484 5160
rect 19892 5108 19944 5160
rect 19984 5108 20036 5160
rect 20812 5244 20864 5296
rect 20720 5176 20772 5228
rect 21088 5244 21140 5296
rect 22284 5244 22336 5296
rect 21272 5176 21324 5228
rect 22468 5176 22520 5228
rect 22652 5219 22704 5228
rect 22652 5185 22661 5219
rect 22661 5185 22695 5219
rect 22695 5185 22704 5219
rect 22652 5176 22704 5185
rect 23388 5176 23440 5228
rect 24032 5176 24084 5228
rect 20812 5108 20864 5160
rect 17776 5040 17828 5049
rect 18880 5040 18932 5092
rect 24952 5176 25004 5228
rect 38016 5219 38068 5228
rect 38016 5185 38025 5219
rect 38025 5185 38059 5219
rect 38059 5185 38068 5219
rect 38016 5176 38068 5185
rect 19892 4972 19944 5024
rect 20628 4972 20680 5024
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 21272 4972 21324 5024
rect 23480 5040 23532 5092
rect 22836 4972 22888 5024
rect 25412 5040 25464 5092
rect 38200 5015 38252 5024
rect 38200 4981 38209 5015
rect 38209 4981 38243 5015
rect 38243 4981 38252 5015
rect 38200 4972 38252 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 3424 4768 3476 4820
rect 4528 4768 4580 4820
rect 5356 4768 5408 4820
rect 8392 4768 8444 4820
rect 10048 4768 10100 4820
rect 10692 4768 10744 4820
rect 12532 4768 12584 4820
rect 3608 4700 3660 4752
rect 4712 4700 4764 4752
rect 1952 4632 2004 4684
rect 3424 4632 3476 4684
rect 3700 4632 3752 4684
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 4712 4564 4764 4616
rect 7012 4564 7064 4616
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 7840 4564 7892 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 12440 4700 12492 4752
rect 12900 4768 12952 4820
rect 13452 4768 13504 4820
rect 14924 4768 14976 4820
rect 17684 4768 17736 4820
rect 18144 4768 18196 4820
rect 18880 4768 18932 4820
rect 8944 4632 8996 4684
rect 10324 4632 10376 4684
rect 11980 4632 12032 4684
rect 14188 4632 14240 4684
rect 14648 4632 14700 4684
rect 3700 4496 3752 4548
rect 5172 4539 5224 4548
rect 5172 4505 5181 4539
rect 5181 4505 5215 4539
rect 5215 4505 5224 4539
rect 5172 4496 5224 4505
rect 5448 4496 5500 4548
rect 9772 4564 9824 4616
rect 10968 4564 11020 4616
rect 14096 4564 14148 4616
rect 19340 4700 19392 4752
rect 19524 4768 19576 4820
rect 19892 4768 19944 4820
rect 20352 4768 20404 4820
rect 20536 4811 20588 4820
rect 20536 4777 20545 4811
rect 20545 4777 20579 4811
rect 20579 4777 20588 4811
rect 20536 4768 20588 4777
rect 21364 4768 21416 4820
rect 23112 4768 23164 4820
rect 23204 4811 23256 4820
rect 23204 4777 23213 4811
rect 23213 4777 23247 4811
rect 23247 4777 23256 4811
rect 23204 4768 23256 4777
rect 22008 4700 22060 4752
rect 24492 4768 24544 4820
rect 28172 4811 28224 4820
rect 16948 4675 17000 4684
rect 16948 4641 16957 4675
rect 16957 4641 16991 4675
rect 16991 4641 17000 4675
rect 16948 4632 17000 4641
rect 17408 4632 17460 4684
rect 17960 4675 18012 4684
rect 16580 4564 16632 4616
rect 17960 4641 17969 4675
rect 17969 4641 18003 4675
rect 18003 4641 18012 4675
rect 17960 4632 18012 4641
rect 18052 4632 18104 4684
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 20168 4632 20220 4684
rect 4988 4428 5040 4480
rect 5264 4428 5316 4480
rect 6920 4428 6972 4480
rect 7932 4428 7984 4480
rect 11428 4496 11480 4548
rect 14280 4496 14332 4548
rect 14556 4539 14608 4548
rect 14556 4505 14565 4539
rect 14565 4505 14599 4539
rect 14599 4505 14608 4539
rect 14556 4496 14608 4505
rect 18604 4564 18656 4616
rect 21272 4632 21324 4684
rect 20352 4564 20404 4616
rect 20536 4496 20588 4548
rect 23388 4632 23440 4684
rect 24860 4700 24912 4752
rect 22468 4607 22520 4616
rect 22468 4573 22477 4607
rect 22477 4573 22511 4607
rect 22511 4573 22520 4607
rect 22468 4564 22520 4573
rect 23112 4607 23164 4616
rect 23112 4573 23121 4607
rect 23121 4573 23155 4607
rect 23155 4573 23164 4607
rect 23112 4564 23164 4573
rect 23296 4564 23348 4616
rect 24768 4632 24820 4684
rect 23572 4564 23624 4616
rect 23848 4607 23900 4616
rect 23848 4573 23857 4607
rect 23857 4573 23891 4607
rect 23891 4573 23900 4607
rect 23848 4564 23900 4573
rect 24492 4564 24544 4616
rect 28172 4777 28181 4811
rect 28181 4777 28215 4811
rect 28215 4777 28224 4811
rect 28172 4768 28224 4777
rect 28264 4768 28316 4820
rect 31392 4768 31444 4820
rect 34060 4768 34112 4820
rect 32312 4700 32364 4752
rect 31392 4607 31444 4616
rect 31392 4573 31401 4607
rect 31401 4573 31435 4607
rect 31435 4573 31444 4607
rect 31392 4564 31444 4573
rect 38292 4607 38344 4616
rect 38292 4573 38301 4607
rect 38301 4573 38335 4607
rect 38335 4573 38344 4607
rect 38292 4564 38344 4573
rect 21088 4496 21140 4548
rect 14924 4428 14976 4480
rect 15936 4428 15988 4480
rect 17316 4428 17368 4480
rect 19892 4428 19944 4480
rect 19984 4428 20036 4480
rect 21364 4428 21416 4480
rect 21640 4428 21692 4480
rect 22008 4428 22060 4480
rect 23112 4428 23164 4480
rect 23664 4496 23716 4548
rect 24584 4428 24636 4480
rect 24768 4428 24820 4480
rect 25044 4471 25096 4480
rect 25044 4437 25053 4471
rect 25053 4437 25087 4471
rect 25087 4437 25096 4471
rect 25044 4428 25096 4437
rect 34428 4428 34480 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2044 4224 2096 4276
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 4896 4224 4948 4276
rect 5080 4224 5132 4276
rect 12900 4224 12952 4276
rect 13820 4224 13872 4276
rect 3424 4199 3476 4208
rect 3424 4165 3433 4199
rect 3433 4165 3467 4199
rect 3467 4165 3476 4199
rect 3424 4156 3476 4165
rect 6460 4156 6512 4208
rect 5724 4088 5776 4140
rect 6184 4088 6236 4140
rect 6828 4156 6880 4208
rect 6920 4156 6972 4208
rect 10876 4156 10928 4208
rect 14004 4156 14056 4208
rect 16856 4224 16908 4276
rect 8300 4088 8352 4140
rect 8852 4088 8904 4140
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 19156 4156 19208 4208
rect 19432 4224 19484 4276
rect 20352 4267 20404 4276
rect 20352 4233 20361 4267
rect 20361 4233 20395 4267
rect 20395 4233 20404 4267
rect 20352 4224 20404 4233
rect 20720 4224 20772 4276
rect 22008 4224 22060 4276
rect 22744 4267 22796 4276
rect 22744 4233 22753 4267
rect 22753 4233 22787 4267
rect 22787 4233 22796 4267
rect 22744 4224 22796 4233
rect 23112 4224 23164 4276
rect 4712 4020 4764 4072
rect 5264 4020 5316 4072
rect 6000 4020 6052 4072
rect 1768 3995 1820 4004
rect 1768 3961 1777 3995
rect 1777 3961 1811 3995
rect 1811 3961 1820 3995
rect 1768 3952 1820 3961
rect 6644 3952 6696 4004
rect 7656 4020 7708 4072
rect 9128 4020 9180 4072
rect 9680 4020 9732 4072
rect 10968 4020 11020 4072
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 13268 4020 13320 4072
rect 14096 4020 14148 4072
rect 14556 4020 14608 4072
rect 13820 3952 13872 4004
rect 6736 3884 6788 3936
rect 9404 3884 9456 3936
rect 11612 3884 11664 3936
rect 11980 3884 12032 3936
rect 12440 3884 12492 3936
rect 17592 4020 17644 4072
rect 17684 4020 17736 4072
rect 19064 4020 19116 4072
rect 16764 3952 16816 4004
rect 19984 4088 20036 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 21180 4020 21232 4072
rect 21272 4020 21324 4072
rect 22192 4088 22244 4140
rect 23756 4088 23808 4140
rect 37188 4156 37240 4208
rect 23020 4020 23072 4072
rect 23204 4020 23256 4072
rect 25780 4088 25832 4140
rect 27344 4131 27396 4140
rect 27344 4097 27353 4131
rect 27353 4097 27387 4131
rect 27387 4097 27396 4131
rect 27344 4088 27396 4097
rect 25136 4020 25188 4072
rect 20812 3952 20864 4004
rect 21732 3952 21784 4004
rect 24768 3952 24820 4004
rect 26884 3952 26936 4004
rect 16304 3884 16356 3936
rect 21640 3884 21692 3936
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 24032 3927 24084 3936
rect 24032 3893 24041 3927
rect 24041 3893 24075 3927
rect 24075 3893 24084 3927
rect 24032 3884 24084 3893
rect 24124 3884 24176 3936
rect 26700 3884 26752 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2504 3680 2556 3732
rect 4068 3680 4120 3732
rect 6092 3680 6144 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 9864 3680 9916 3732
rect 11980 3680 12032 3732
rect 12256 3680 12308 3732
rect 13176 3680 13228 3732
rect 14556 3680 14608 3732
rect 19892 3680 19944 3732
rect 20168 3723 20220 3732
rect 20168 3689 20177 3723
rect 20177 3689 20211 3723
rect 20211 3689 20220 3723
rect 20168 3680 20220 3689
rect 20628 3680 20680 3732
rect 24676 3680 24728 3732
rect 25872 3680 25924 3732
rect 4344 3612 4396 3664
rect 7012 3612 7064 3664
rect 8576 3612 8628 3664
rect 11612 3612 11664 3664
rect 13544 3612 13596 3664
rect 14280 3612 14332 3664
rect 18972 3612 19024 3664
rect 4344 3476 4396 3528
rect 6736 3544 6788 3596
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 4436 3340 4488 3392
rect 6828 3476 6880 3528
rect 7656 3476 7708 3528
rect 8300 3476 8352 3528
rect 9588 3476 9640 3528
rect 11796 3544 11848 3596
rect 12348 3587 12400 3596
rect 12348 3553 12357 3587
rect 12357 3553 12391 3587
rect 12391 3553 12400 3587
rect 12348 3544 12400 3553
rect 16120 3544 16172 3596
rect 16948 3544 17000 3596
rect 20076 3612 20128 3664
rect 20352 3612 20404 3664
rect 22100 3655 22152 3664
rect 22100 3621 22109 3655
rect 22109 3621 22143 3655
rect 22143 3621 22152 3655
rect 22100 3612 22152 3621
rect 37740 3680 37792 3732
rect 19340 3544 19392 3596
rect 20536 3544 20588 3596
rect 20812 3587 20864 3596
rect 20812 3553 20821 3587
rect 20821 3553 20855 3587
rect 20855 3553 20864 3587
rect 20812 3544 20864 3553
rect 21916 3544 21968 3596
rect 11980 3476 12032 3528
rect 16764 3519 16816 3528
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 17040 3476 17092 3528
rect 18696 3476 18748 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 4804 3451 4856 3460
rect 4804 3417 4813 3451
rect 4813 3417 4847 3451
rect 4847 3417 4856 3451
rect 4804 3408 4856 3417
rect 4896 3340 4948 3392
rect 6644 3408 6696 3460
rect 12164 3408 12216 3460
rect 14280 3408 14332 3460
rect 7012 3340 7064 3392
rect 8668 3340 8720 3392
rect 11244 3340 11296 3392
rect 13360 3340 13412 3392
rect 14556 3451 14608 3460
rect 14556 3417 14565 3451
rect 14565 3417 14599 3451
rect 14599 3417 14608 3451
rect 14556 3408 14608 3417
rect 15200 3408 15252 3460
rect 14740 3340 14792 3392
rect 15844 3408 15896 3460
rect 17776 3451 17828 3460
rect 17776 3417 17785 3451
rect 17785 3417 17819 3451
rect 17819 3417 17828 3451
rect 17776 3408 17828 3417
rect 17684 3340 17736 3392
rect 19708 3408 19760 3460
rect 20076 3340 20128 3392
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 21456 3476 21508 3528
rect 20536 3408 20588 3460
rect 21088 3408 21140 3460
rect 25044 3544 25096 3596
rect 22468 3476 22520 3528
rect 24216 3476 24268 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 25136 3476 25188 3528
rect 25780 3476 25832 3528
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 27436 3408 27488 3460
rect 37924 3476 37976 3528
rect 22192 3340 22244 3392
rect 23480 3340 23532 3392
rect 24860 3340 24912 3392
rect 26608 3383 26660 3392
rect 26608 3349 26617 3383
rect 26617 3349 26651 3383
rect 26651 3349 26660 3383
rect 26608 3340 26660 3349
rect 27160 3383 27212 3392
rect 27160 3349 27169 3383
rect 27169 3349 27203 3383
rect 27203 3349 27212 3383
rect 27160 3340 27212 3349
rect 27804 3383 27856 3392
rect 27804 3349 27813 3383
rect 27813 3349 27847 3383
rect 27847 3349 27856 3383
rect 27804 3340 27856 3349
rect 38016 3340 38068 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4436 3136 4488 3188
rect 5448 3136 5500 3188
rect 7564 3136 7616 3188
rect 8116 3136 8168 3188
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 12808 3136 12860 3188
rect 13452 3136 13504 3188
rect 2412 3068 2464 3120
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 5540 3068 5592 3120
rect 6644 3068 6696 3120
rect 7196 3068 7248 3120
rect 5172 3043 5224 3052
rect 20 2864 72 2916
rect 664 2796 716 2848
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 6552 3000 6604 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 5632 2932 5684 2984
rect 6460 2932 6512 2984
rect 4436 2864 4488 2916
rect 7196 2864 7248 2916
rect 7840 3000 7892 3052
rect 8208 3000 8260 3052
rect 7932 2932 7984 2984
rect 10232 3000 10284 3052
rect 10692 3000 10744 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 11060 2932 11112 2984
rect 11428 2932 11480 2984
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 13728 2932 13780 2984
rect 5724 2796 5776 2848
rect 6368 2796 6420 2848
rect 11244 2864 11296 2916
rect 12716 2796 12768 2848
rect 15108 3136 15160 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 16028 3179 16080 3188
rect 16028 3145 16037 3179
rect 16037 3145 16071 3179
rect 16071 3145 16080 3179
rect 16028 3136 16080 3145
rect 16396 3136 16448 3188
rect 18420 3179 18472 3188
rect 14924 3068 14976 3120
rect 16488 3068 16540 3120
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 18512 3136 18564 3188
rect 19156 3136 19208 3188
rect 20812 3136 20864 3188
rect 21364 3136 21416 3188
rect 30748 3136 30800 3188
rect 16764 3000 16816 3052
rect 18328 3043 18380 3052
rect 18328 3009 18337 3043
rect 18337 3009 18371 3043
rect 18371 3009 18380 3043
rect 18328 3000 18380 3009
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 19616 3041 19668 3052
rect 19616 3007 19633 3041
rect 19633 3007 19667 3041
rect 19667 3007 19668 3041
rect 19616 3000 19668 3007
rect 20168 3000 20220 3052
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 22376 3068 22428 3120
rect 24676 3068 24728 3120
rect 25504 3111 25556 3120
rect 25504 3077 25513 3111
rect 25513 3077 25547 3111
rect 25547 3077 25556 3111
rect 25504 3068 25556 3077
rect 22652 3043 22704 3052
rect 18236 2932 18288 2984
rect 19340 2932 19392 2984
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 22284 2932 22336 2984
rect 22928 2932 22980 2984
rect 15292 2796 15344 2848
rect 15660 2796 15712 2848
rect 16120 2796 16172 2848
rect 17316 2864 17368 2916
rect 20536 2864 20588 2916
rect 25320 3000 25372 3052
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 25688 3000 25740 3052
rect 27988 3043 28040 3052
rect 24216 2932 24268 2984
rect 27436 2932 27488 2984
rect 21824 2796 21876 2848
rect 21916 2796 21968 2848
rect 24584 2864 24636 2916
rect 27988 3009 27997 3043
rect 27997 3009 28031 3043
rect 28031 3009 28040 3043
rect 27988 3000 28040 3009
rect 37740 3043 37792 3052
rect 37464 2975 37516 2984
rect 37464 2941 37473 2975
rect 37473 2941 37507 2975
rect 37507 2941 37516 2975
rect 37464 2932 37516 2941
rect 37740 3009 37749 3043
rect 37749 3009 37783 3043
rect 37783 3009 37792 3043
rect 37740 3000 37792 3009
rect 39304 2932 39356 2984
rect 22744 2839 22796 2848
rect 22744 2805 22753 2839
rect 22753 2805 22787 2839
rect 22787 2805 22796 2839
rect 22744 2796 22796 2805
rect 23296 2839 23348 2848
rect 23296 2805 23305 2839
rect 23305 2805 23339 2839
rect 23339 2805 23348 2839
rect 23296 2796 23348 2805
rect 26056 2839 26108 2848
rect 26056 2805 26065 2839
rect 26065 2805 26099 2839
rect 26099 2805 26108 2839
rect 26056 2796 26108 2805
rect 27252 2839 27304 2848
rect 27252 2805 27261 2839
rect 27261 2805 27295 2839
rect 27295 2805 27304 2839
rect 27252 2796 27304 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 7012 2592 7064 2644
rect 5448 2524 5500 2576
rect 9956 2592 10008 2644
rect 10140 2592 10192 2644
rect 12624 2592 12676 2644
rect 13728 2635 13780 2644
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 16120 2635 16172 2644
rect 16120 2601 16129 2635
rect 16129 2601 16163 2635
rect 16163 2601 16172 2635
rect 16120 2592 16172 2601
rect 16488 2592 16540 2644
rect 17500 2592 17552 2644
rect 20352 2592 20404 2644
rect 22652 2592 22704 2644
rect 24308 2592 24360 2644
rect 25320 2592 25372 2644
rect 28448 2635 28500 2644
rect 28448 2601 28457 2635
rect 28457 2601 28491 2635
rect 28491 2601 28500 2635
rect 28448 2592 28500 2601
rect 30472 2635 30524 2644
rect 30472 2601 30481 2635
rect 30481 2601 30515 2635
rect 30515 2601 30524 2635
rect 30472 2592 30524 2601
rect 32312 2635 32364 2644
rect 32312 2601 32321 2635
rect 32321 2601 32355 2635
rect 32355 2601 32364 2635
rect 32312 2592 32364 2601
rect 33140 2635 33192 2644
rect 33140 2601 33149 2635
rect 33149 2601 33183 2635
rect 33183 2601 33192 2635
rect 33140 2592 33192 2601
rect 8300 2524 8352 2576
rect 9220 2456 9272 2508
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 3884 2388 3936 2440
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 7196 2388 7248 2440
rect 8208 2388 8260 2440
rect 4620 2320 4672 2372
rect 8484 2388 8536 2440
rect 15844 2524 15896 2576
rect 11704 2456 11756 2508
rect 13544 2456 13596 2508
rect 15384 2431 15436 2440
rect 15384 2397 15393 2431
rect 15393 2397 15427 2431
rect 15427 2397 15436 2431
rect 15384 2388 15436 2397
rect 15936 2388 15988 2440
rect 16304 2388 16356 2440
rect 16948 2388 17000 2440
rect 19432 2524 19484 2576
rect 19248 2456 19300 2508
rect 23480 2524 23532 2576
rect 21824 2456 21876 2508
rect 20076 2431 20128 2440
rect 8576 2320 8628 2372
rect 9956 2320 10008 2372
rect 10508 2320 10560 2372
rect 17960 2320 18012 2372
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20628 2388 20680 2440
rect 21916 2388 21968 2440
rect 31116 2456 31168 2508
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 23848 2388 23900 2440
rect 25596 2388 25648 2440
rect 25964 2431 26016 2440
rect 25964 2397 25973 2431
rect 25973 2397 26007 2431
rect 26007 2397 26016 2431
rect 25964 2388 26016 2397
rect 27068 2388 27120 2440
rect 28356 2388 28408 2440
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 30288 2388 30340 2440
rect 31576 2388 31628 2440
rect 33692 2431 33744 2440
rect 33692 2397 33701 2431
rect 33701 2397 33735 2431
rect 33735 2397 33744 2431
rect 33692 2388 33744 2397
rect 34428 2388 34480 2440
rect 36728 2388 36780 2440
rect 37740 2431 37792 2440
rect 37740 2397 37749 2431
rect 37749 2397 37783 2431
rect 37783 2397 37792 2431
rect 37740 2388 37792 2397
rect 23296 2320 23348 2372
rect 32864 2320 32916 2372
rect 1952 2252 2004 2304
rect 3240 2252 3292 2304
rect 5172 2252 5224 2304
rect 6460 2252 6512 2304
rect 13084 2252 13136 2304
rect 15476 2295 15528 2304
rect 15476 2261 15485 2295
rect 15485 2261 15519 2295
rect 15519 2261 15528 2295
rect 15476 2252 15528 2261
rect 18052 2252 18104 2304
rect 20996 2252 21048 2304
rect 22560 2252 22612 2304
rect 23388 2295 23440 2304
rect 23388 2261 23397 2295
rect 23397 2261 23431 2295
rect 23431 2261 23440 2295
rect 23388 2252 23440 2261
rect 25136 2252 25188 2304
rect 25780 2252 25832 2304
rect 29644 2252 29696 2304
rect 33508 2252 33560 2304
rect 34796 2252 34848 2304
rect 36084 2252 36136 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 10876 2048 10928 2100
rect 27252 2048 27304 2100
rect 3608 1980 3660 2032
rect 15476 1980 15528 2032
rect 17960 1980 18012 2032
rect 24860 1980 24912 2032
rect 10784 1912 10836 1964
rect 9036 1844 9088 1896
rect 19248 1844 19300 1896
rect 20076 1912 20128 1964
rect 26700 1912 26752 1964
rect 24124 1844 24176 1896
rect 8576 1776 8628 1828
rect 15384 1776 15436 1828
rect 13728 1708 13780 1760
rect 22192 1708 22244 1760
rect 22284 1708 22336 1760
rect 37740 1776 37792 1828
rect 16120 1640 16172 1692
rect 17316 1640 17368 1692
rect 17408 1640 17460 1692
rect 23572 1640 23624 1692
rect 13820 1572 13872 1624
rect 21548 1572 21600 1624
rect 20536 1300 20588 1352
rect 25688 1300 25740 1352
rect 14832 1232 14884 1284
rect 24768 1232 24820 1284
rect 4988 1164 5040 1216
rect 21272 1164 21324 1216
rect 10876 144 10928 196
rect 24952 144 25004 196
rect 11704 76 11756 128
rect 27988 76 28040 128
rect 7196 8 7248 60
rect 27344 8 27396 60
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14186 39200 14242 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 17406 39200 17462 39800
rect 18694 39200 18750 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25134 39200 25190 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28354 39200 28410 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 32 36786 60 39200
rect 1320 36854 1348 39200
rect 1582 38856 1638 38865
rect 1582 38791 1638 38800
rect 1596 37330 1624 38791
rect 1766 38176 1822 38185
rect 1766 38111 1822 38120
rect 1584 37324 1636 37330
rect 1584 37266 1636 37272
rect 1308 36848 1360 36854
rect 1308 36790 1360 36796
rect 20 36780 72 36786
rect 20 36722 72 36728
rect 1780 36378 1808 38111
rect 2608 37210 2636 39200
rect 3252 37262 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 37726
rect 5828 37262 5856 39200
rect 6472 37262 6500 39200
rect 2872 37256 2924 37262
rect 2608 37182 2820 37210
rect 2872 37198 2924 37204
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 5540 37256 5592 37262
rect 5540 37198 5592 37204
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 2792 37126 2820 37182
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 1860 36712 1912 36718
rect 1860 36654 1912 36660
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1596 36009 1624 36110
rect 1582 36000 1638 36009
rect 1582 35935 1638 35944
rect 1768 35488 1820 35494
rect 1766 35456 1768 35465
rect 1820 35456 1822 35465
rect 1766 35391 1822 35400
rect 1768 35080 1820 35086
rect 1768 35022 1820 35028
rect 1780 34785 1808 35022
rect 1766 34776 1822 34785
rect 1766 34711 1822 34720
rect 1766 33416 1822 33425
rect 1766 33351 1768 33360
rect 1820 33351 1822 33360
rect 1768 33322 1820 33328
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1596 32065 1624 32302
rect 1582 32056 1638 32065
rect 1582 31991 1638 32000
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1780 31385 1808 31622
rect 1766 31376 1822 31385
rect 1766 31311 1822 31320
rect 1872 30666 1900 36654
rect 2792 36174 2820 36751
rect 2780 36168 2832 36174
rect 2780 36110 2832 36116
rect 1860 30660 1912 30666
rect 1860 30602 1912 30608
rect 1768 30048 1820 30054
rect 1766 30016 1768 30025
rect 1820 30016 1822 30025
rect 1766 29951 1822 29960
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1780 28665 1808 29106
rect 2688 29028 2740 29034
rect 2688 28970 2740 28976
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 26625 1440 28018
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 1768 27328 1820 27334
rect 1766 27296 1768 27305
rect 1820 27296 1822 27305
rect 1766 27231 1822 27240
rect 1860 26988 1912 26994
rect 1860 26930 1912 26936
rect 2320 26988 2372 26994
rect 2320 26930 2372 26936
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1398 26616 1454 26625
rect 1398 26551 1454 26560
rect 1124 25900 1176 25906
rect 1124 25842 1176 25848
rect 1032 25220 1084 25226
rect 1032 25162 1084 25168
rect 940 24404 992 24410
rect 940 24346 992 24352
rect 952 10742 980 24346
rect 1044 11082 1072 25162
rect 1136 12209 1164 25842
rect 1216 25832 1268 25838
rect 1216 25774 1268 25780
rect 1122 12200 1178 12209
rect 1122 12135 1178 12144
rect 1228 11694 1256 25774
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1492 24200 1544 24206
rect 1492 24142 1544 24148
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1308 23588 1360 23594
rect 1308 23530 1360 23536
rect 1320 20602 1348 23530
rect 1308 20596 1360 20602
rect 1308 20538 1360 20544
rect 1216 11688 1268 11694
rect 1216 11630 1268 11636
rect 1032 11076 1084 11082
rect 1032 11018 1084 11024
rect 1308 11076 1360 11082
rect 1308 11018 1360 11024
rect 940 10736 992 10742
rect 940 10678 992 10684
rect 952 7954 980 10678
rect 1320 8362 1348 11018
rect 1412 8634 1440 23666
rect 1504 16998 1532 24142
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21865 1624 21966
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 1688 20534 1716 26726
rect 1872 26625 1900 26930
rect 2332 26897 2360 26930
rect 2318 26888 2374 26897
rect 2318 26823 2374 26832
rect 1858 26616 1914 26625
rect 1858 26551 1914 26560
rect 2228 26376 2280 26382
rect 2228 26318 2280 26324
rect 1860 25696 1912 25702
rect 1860 25638 1912 25644
rect 1768 23044 1820 23050
rect 1768 22986 1820 22992
rect 1676 20528 1728 20534
rect 1676 20470 1728 20476
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1596 18222 1624 18702
rect 1584 18216 1636 18222
rect 1636 18176 1716 18204
rect 1584 18158 1636 18164
rect 1688 17746 1716 18176
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1584 17128 1636 17134
rect 1688 17116 1716 17682
rect 1636 17088 1716 17116
rect 1584 17070 1636 17076
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16794 1532 16934
rect 1492 16788 1544 16794
rect 1492 16730 1544 16736
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1596 16640 1624 16730
rect 1688 16658 1716 17088
rect 1504 16612 1624 16640
rect 1676 16652 1728 16658
rect 1504 8974 1532 16612
rect 1676 16594 1728 16600
rect 1688 16114 1716 16594
rect 1780 16574 1808 22986
rect 1872 21622 1900 25638
rect 1952 24880 2004 24886
rect 1952 24822 2004 24828
rect 1860 21616 1912 21622
rect 1860 21558 1912 21564
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 1872 19854 1900 21082
rect 1964 20534 1992 24822
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 2056 23526 2084 24550
rect 2136 23656 2188 23662
rect 2134 23624 2136 23633
rect 2188 23624 2190 23633
rect 2134 23559 2190 23568
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2148 21146 2176 22510
rect 2136 21140 2188 21146
rect 2136 21082 2188 21088
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 1952 20528 2004 20534
rect 1952 20470 2004 20476
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1858 17368 1914 17377
rect 1858 17303 1914 17312
rect 1872 17270 1900 17303
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 1964 17134 1992 17546
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2056 16794 2084 20538
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 1780 16546 1900 16574
rect 1676 16108 1728 16114
rect 1596 16068 1676 16096
rect 1596 15570 1624 16068
rect 1676 16050 1728 16056
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1596 15026 1624 15506
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 14482 1624 14962
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 12782 1624 13330
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1596 12306 1624 12718
rect 1872 12434 1900 16546
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1688 12406 1900 12434
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1596 11762 1624 12242
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 11218 1624 11698
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1308 8356 1360 8362
rect 1308 8298 1360 8304
rect 1688 8090 1716 12406
rect 1858 11928 1914 11937
rect 1964 11898 1992 15302
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1858 11863 1914 11872
rect 1952 11892 2004 11898
rect 1872 11830 1900 11863
rect 1952 11834 2004 11840
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 10810 1808 10950
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1964 9994 1992 11630
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1780 8838 1808 8871
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 940 7948 992 7954
rect 940 7890 992 7896
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7585 1624 7822
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 20 2916 72 2922
rect 20 2858 72 2864
rect 32 800 60 2858
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 676 800 704 2790
rect 18 200 74 800
rect 662 200 718 800
rect 1412 785 1440 7346
rect 2056 7002 2084 12582
rect 2148 9110 2176 19382
rect 2240 16574 2268 26318
rect 2320 26308 2372 26314
rect 2320 26250 2372 26256
rect 2332 20874 2360 26250
rect 2320 20868 2372 20874
rect 2320 20810 2372 20816
rect 2424 18034 2452 27406
rect 2504 27328 2556 27334
rect 2504 27270 2556 27276
rect 2516 24886 2544 27270
rect 2596 26784 2648 26790
rect 2596 26726 2648 26732
rect 2504 24880 2556 24886
rect 2504 24822 2556 24828
rect 2504 24200 2556 24206
rect 2502 24168 2504 24177
rect 2556 24168 2558 24177
rect 2502 24103 2558 24112
rect 2504 24064 2556 24070
rect 2504 24006 2556 24012
rect 2516 22166 2544 24006
rect 2608 22982 2636 26726
rect 2700 26466 2728 28970
rect 2884 28490 2912 37198
rect 3976 37120 4028 37126
rect 3976 37062 4028 37068
rect 3988 29714 4016 37062
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4620 35692 4672 35698
rect 4620 35634 4672 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 34944 4120 34950
rect 4068 34886 4120 34892
rect 4080 30734 4108 34886
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 32026 4660 35634
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30728 4120 30734
rect 4068 30670 4120 30676
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3976 29708 4028 29714
rect 3976 29650 4028 29656
rect 4632 29306 4660 31758
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 4620 29300 4672 29306
rect 4620 29242 4672 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 2872 28484 2924 28490
rect 2872 28426 2924 28432
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3240 26784 3292 26790
rect 3240 26726 3292 26732
rect 2700 26438 2820 26466
rect 2688 26376 2740 26382
rect 2686 26344 2688 26353
rect 2740 26344 2742 26353
rect 2686 26279 2742 26288
rect 2792 26234 2820 26438
rect 3252 26353 3280 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4068 26512 4120 26518
rect 4068 26454 4120 26460
rect 3238 26344 3294 26353
rect 2964 26308 3016 26314
rect 3238 26279 3294 26288
rect 2964 26250 3016 26256
rect 2700 26206 2820 26234
rect 2700 24818 2728 26206
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2504 22160 2556 22166
rect 2504 22102 2556 22108
rect 2594 20632 2650 20641
rect 2594 20567 2650 20576
rect 2608 20534 2636 20567
rect 2596 20528 2648 20534
rect 2596 20470 2648 20476
rect 2504 19780 2556 19786
rect 2504 19722 2556 19728
rect 2332 18006 2452 18034
rect 2332 17490 2360 18006
rect 2332 17462 2452 17490
rect 2240 16546 2360 16574
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2240 13705 2268 13874
rect 2226 13696 2282 13705
rect 2226 13631 2282 13640
rect 2332 11558 2360 16546
rect 2424 14958 2452 17462
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2318 10840 2374 10849
rect 2516 10810 2544 19722
rect 2608 19446 2636 20470
rect 2596 19440 2648 19446
rect 2596 19382 2648 19388
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2608 15366 2636 17274
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2608 14278 2636 14894
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2700 13870 2728 23462
rect 2792 22710 2820 24550
rect 2780 22704 2832 22710
rect 2780 22646 2832 22652
rect 2884 22556 2912 25774
rect 2976 23186 3004 26250
rect 3792 25696 3844 25702
rect 3976 25696 4028 25702
rect 3792 25638 3844 25644
rect 3974 25664 3976 25673
rect 4028 25664 4030 25673
rect 3240 25152 3292 25158
rect 3240 25094 3292 25100
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 3068 23594 3096 24550
rect 3148 24064 3200 24070
rect 3148 24006 3200 24012
rect 3056 23588 3108 23594
rect 3056 23530 3108 23536
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 3056 23112 3108 23118
rect 3056 23054 3108 23060
rect 2792 22528 2912 22556
rect 2792 21078 2820 22528
rect 3068 22386 3096 23054
rect 2884 22358 3096 22386
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2792 16046 2820 18362
rect 2884 18154 2912 22358
rect 3160 22080 3188 24006
rect 3252 22778 3280 25094
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3332 24064 3384 24070
rect 3332 24006 3384 24012
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3252 22234 3280 22374
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3240 22092 3292 22098
rect 3160 22052 3240 22080
rect 3240 22034 3292 22040
rect 3238 21992 3294 22001
rect 2964 21956 3016 21962
rect 3238 21927 3294 21936
rect 2964 21898 3016 21904
rect 2976 20505 3004 21898
rect 3252 21894 3280 21927
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3252 21146 3280 21626
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 2962 20496 3018 20505
rect 2962 20431 3018 20440
rect 3344 20398 3372 24006
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 2872 18148 2924 18154
rect 2872 18090 2924 18096
rect 2884 16454 2912 18090
rect 3056 17808 3108 17814
rect 3056 17750 3108 17756
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2792 14074 2820 15671
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2976 13530 3004 17002
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2870 11656 2926 11665
rect 2870 11591 2926 11600
rect 2318 10775 2320 10784
rect 2372 10775 2374 10784
rect 2504 10804 2556 10810
rect 2320 10746 2372 10752
rect 2504 10746 2556 10752
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2240 8430 2268 9318
rect 2516 9058 2544 9454
rect 2608 9382 2636 10066
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2594 9208 2650 9217
rect 2594 9143 2596 9152
rect 2648 9143 2650 9152
rect 2688 9172 2740 9178
rect 2596 9114 2648 9120
rect 2688 9114 2740 9120
rect 2700 9058 2728 9114
rect 2516 9030 2728 9058
rect 2792 8974 2820 10231
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 7410 2268 8366
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 5778 1624 6734
rect 1950 6352 2006 6361
rect 1950 6287 1952 6296
rect 2004 6287 2006 6296
rect 1952 6258 2004 6264
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 2056 5166 2084 5714
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1952 4684 2004 4690
rect 2056 4672 2084 5102
rect 2004 4644 2084 4672
rect 1952 4626 2004 4632
rect 2056 4282 2084 4644
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 1766 4176 1822 4185
rect 1584 4140 1636 4146
rect 1766 4111 1822 4120
rect 1584 4082 1636 4088
rect 1596 3369 1624 4082
rect 1780 4010 1808 4111
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 1768 3392 1820 3398
rect 1582 3360 1638 3369
rect 1768 3334 1820 3340
rect 1582 3295 1638 3304
rect 1780 2145 1808 3334
rect 2332 3058 2360 6054
rect 2424 3126 2452 6054
rect 2516 3738 2544 8910
rect 2884 8634 2912 11591
rect 3068 10674 3096 17750
rect 3160 16266 3188 18634
rect 3252 18465 3280 19314
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18834 3372 19110
rect 3436 18970 3464 24754
rect 3712 24410 3740 24754
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3804 24188 3832 25638
rect 3974 25599 4030 25608
rect 3976 25288 4028 25294
rect 3976 25230 4028 25236
rect 3988 24993 4016 25230
rect 3974 24984 4030 24993
rect 3974 24919 4030 24928
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3896 24342 3924 24550
rect 3884 24336 3936 24342
rect 3884 24278 3936 24284
rect 3804 24160 3924 24188
rect 3608 24132 3660 24138
rect 3608 24074 3660 24080
rect 3620 23866 3648 24074
rect 3608 23860 3660 23866
rect 3608 23802 3660 23808
rect 3608 23656 3660 23662
rect 3608 23598 3660 23604
rect 3516 23248 3568 23254
rect 3514 23216 3516 23225
rect 3568 23216 3570 23225
rect 3514 23151 3570 23160
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3528 22710 3556 22918
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3620 22250 3648 23598
rect 3698 23080 3754 23089
rect 3698 23015 3754 23024
rect 3792 23044 3844 23050
rect 3528 22222 3648 22250
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3330 18592 3386 18601
rect 3330 18527 3386 18536
rect 3238 18456 3294 18465
rect 3344 18426 3372 18527
rect 3238 18391 3294 18400
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3436 18222 3464 18906
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3330 17912 3386 17921
rect 3330 17847 3386 17856
rect 3160 16238 3280 16266
rect 3252 15586 3280 16238
rect 3344 16182 3372 17847
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3160 15558 3280 15586
rect 3424 15564 3476 15570
rect 3160 12442 3188 15558
rect 3424 15506 3476 15512
rect 3436 15337 3464 15506
rect 3422 15328 3478 15337
rect 3422 15263 3478 15272
rect 3332 14952 3384 14958
rect 3330 14920 3332 14929
rect 3384 14920 3386 14929
rect 3330 14855 3386 14864
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3252 12345 3280 13670
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3344 12986 3372 13466
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3332 12776 3384 12782
rect 3330 12744 3332 12753
rect 3384 12744 3386 12753
rect 3330 12679 3386 12688
rect 3332 12436 3384 12442
rect 3528 12434 3556 22222
rect 3608 22092 3660 22098
rect 3608 22034 3660 22040
rect 3620 21486 3648 22034
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3712 19718 3740 23015
rect 3792 22986 3844 22992
rect 3804 22506 3832 22986
rect 3896 22545 3924 24160
rect 3976 23588 4028 23594
rect 3976 23530 4028 23536
rect 3882 22536 3938 22545
rect 3792 22500 3844 22506
rect 3882 22471 3938 22480
rect 3792 22442 3844 22448
rect 3988 22420 4016 23530
rect 4080 23118 4108 26454
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 4540 24818 4568 25230
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4528 24812 4580 24818
rect 4528 24754 4580 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4344 24268 4396 24274
rect 4344 24210 4396 24216
rect 4356 23526 4384 24210
rect 4632 23798 4660 25094
rect 4724 24206 4752 25638
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4712 24064 4764 24070
rect 4712 24006 4764 24012
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4344 23520 4396 23526
rect 4344 23462 4396 23468
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 3896 22392 4016 22420
rect 4068 22432 4120 22438
rect 3896 22386 3924 22392
rect 3804 22358 3924 22386
rect 4068 22374 4120 22380
rect 3804 21486 3832 22358
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21690 4016 21966
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 3882 21584 3938 21593
rect 3882 21519 3938 21528
rect 3792 21480 3844 21486
rect 3792 21422 3844 21428
rect 3790 20768 3846 20777
rect 3790 20703 3846 20712
rect 3700 19712 3752 19718
rect 3606 19680 3662 19689
rect 3700 19654 3752 19660
rect 3606 19615 3662 19624
rect 3620 17134 3648 19615
rect 3698 19544 3754 19553
rect 3698 19479 3700 19488
rect 3752 19479 3754 19488
rect 3700 19450 3752 19456
rect 3804 18714 3832 20703
rect 3712 18686 3832 18714
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3620 16969 3648 17070
rect 3606 16960 3662 16969
rect 3606 16895 3662 16904
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3620 15706 3648 16594
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3620 15162 3648 15642
rect 3712 15450 3740 18686
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3804 17814 3832 18566
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 3790 17504 3846 17513
rect 3790 17439 3846 17448
rect 3804 17202 3832 17439
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3896 16590 3924 21519
rect 3974 20632 4030 20641
rect 3974 20567 4030 20576
rect 3988 20534 4016 20567
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18766 4016 19314
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3988 17882 4016 18702
rect 4080 18426 4108 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22094 4660 23462
rect 4540 22066 4660 22094
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4172 21622 4200 21830
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4264 21457 4292 21966
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 4448 21729 4476 21898
rect 4434 21720 4490 21729
rect 4434 21655 4490 21664
rect 4250 21448 4306 21457
rect 4250 21383 4306 21392
rect 4540 21350 4568 22066
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21026 4660 21966
rect 4724 21894 4752 24006
rect 4816 23254 4844 26318
rect 4896 25900 4948 25906
rect 4896 25842 4948 25848
rect 4908 23905 4936 25842
rect 4988 24608 5040 24614
rect 4988 24550 5040 24556
rect 5000 24206 5028 24550
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 4988 24064 5040 24070
rect 4986 24032 4988 24041
rect 5040 24032 5042 24041
rect 4986 23967 5042 23976
rect 4894 23896 4950 23905
rect 4894 23831 4950 23840
rect 5184 23798 5212 27814
rect 5264 27396 5316 27402
rect 5264 27338 5316 27344
rect 5276 25498 5304 27338
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5356 25288 5408 25294
rect 5356 25230 5408 25236
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5172 23792 5224 23798
rect 5172 23734 5224 23740
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 4804 23248 4856 23254
rect 4804 23190 4856 23196
rect 4894 22536 4950 22545
rect 4894 22471 4950 22480
rect 4804 22160 4856 22166
rect 4804 22102 4856 22108
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4712 21412 4764 21418
rect 4712 21354 4764 21360
rect 4724 21078 4752 21354
rect 4448 20998 4660 21026
rect 4712 21072 4764 21078
rect 4712 21014 4764 21020
rect 4448 20602 4476 20998
rect 4526 20904 4582 20913
rect 4526 20839 4528 20848
rect 4580 20839 4582 20848
rect 4528 20810 4580 20816
rect 4724 20754 4752 21014
rect 4816 20874 4844 22102
rect 4908 21690 4936 22471
rect 5092 22094 5120 23666
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5000 22066 5120 22094
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 4804 20868 4856 20874
rect 4804 20810 4856 20816
rect 4896 20800 4948 20806
rect 4724 20726 4844 20754
rect 4896 20742 4948 20748
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4712 20324 4764 20330
rect 4712 20266 4764 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4724 19922 4752 20266
rect 4816 20058 4844 20726
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4712 19916 4764 19922
rect 4712 19858 4764 19864
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4356 19553 4384 19790
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4342 19544 4398 19553
rect 4342 19479 4398 19488
rect 4724 19310 4752 19654
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3974 17776 4030 17785
rect 3974 17711 4030 17720
rect 3988 17066 4016 17711
rect 4080 17270 4108 17818
rect 4526 17640 4582 17649
rect 4252 17604 4304 17610
rect 4526 17575 4582 17584
rect 4252 17546 4304 17552
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4264 17082 4292 17546
rect 4540 17270 4568 17575
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 4632 17134 4660 18294
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 4080 17054 4292 17082
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4080 16708 4108 17054
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4160 16720 4212 16726
rect 4080 16680 4160 16708
rect 4160 16662 4212 16668
rect 4632 16658 4660 17070
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 3790 16280 3846 16289
rect 3790 16215 3792 16224
rect 3844 16215 3846 16224
rect 3792 16186 3844 16192
rect 3712 15422 3924 15450
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3332 12378 3384 12384
rect 3436 12406 3556 12434
rect 3238 12336 3294 12345
rect 3238 12271 3294 12280
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2976 8566 3004 10202
rect 3252 9081 3280 12038
rect 3344 10810 3372 12378
rect 3436 12102 3464 12406
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3436 10742 3464 12038
rect 3528 11694 3556 12038
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3620 11694 3648 11834
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11218 3556 11494
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3528 9994 3556 11154
rect 3620 10577 3648 11630
rect 3606 10568 3662 10577
rect 3606 10503 3662 10512
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3238 9072 3294 9081
rect 3238 9007 3294 9016
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2870 7984 2926 7993
rect 2870 7919 2926 7928
rect 2884 7886 2912 7919
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3344 5574 3372 6802
rect 3436 5914 3464 9318
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 2688 5160 2740 5166
rect 2686 5128 2688 5137
rect 2740 5128 2742 5137
rect 2686 5063 2742 5072
rect 3436 4826 3464 5510
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3436 4214 3464 4626
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 3528 2774 3556 9590
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3620 6633 3648 9046
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3606 6624 3662 6633
rect 3606 6559 3662 6568
rect 3620 4758 3648 6559
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3712 4690 3740 8298
rect 3804 7954 3832 10474
rect 3896 9382 3924 15422
rect 3988 13326 4016 16458
rect 4264 16114 4292 16458
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 16594
rect 4724 16522 4752 17682
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4172 15094 4200 15370
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 13954 4292 14418
rect 4172 13938 4292 13954
rect 4160 13932 4292 13938
rect 4212 13926 4292 13932
rect 4160 13874 4212 13880
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13394 4660 13670
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12073 4016 13126
rect 4068 12912 4120 12918
rect 4066 12880 4068 12889
rect 4120 12880 4122 12889
rect 4066 12815 4122 12824
rect 4172 12782 4200 13262
rect 4632 13258 4660 13330
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4160 12776 4212 12782
rect 4080 12724 4160 12730
rect 4080 12718 4212 12724
rect 4080 12702 4200 12718
rect 4080 12442 4108 12702
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4264 12209 4292 12242
rect 4250 12200 4306 12209
rect 4160 12164 4212 12170
rect 4250 12135 4252 12144
rect 4160 12106 4212 12112
rect 4304 12135 4306 12144
rect 4252 12106 4304 12112
rect 3974 12064 4030 12073
rect 3974 11999 4030 12008
rect 4172 11898 4200 12106
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4632 11830 4660 13194
rect 4724 12442 4752 14758
rect 4816 14550 4844 19858
rect 4908 17354 4936 20742
rect 5000 20602 5028 22066
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5092 21865 5120 21966
rect 5078 21856 5134 21865
rect 5078 21791 5134 21800
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 5000 17542 5028 19246
rect 5092 17610 5120 21626
rect 5184 19786 5212 23462
rect 5172 19780 5224 19786
rect 5172 19722 5224 19728
rect 5276 19446 5304 24550
rect 5368 23089 5396 25230
rect 5460 23866 5488 30194
rect 5552 24818 5580 37198
rect 7760 37126 7788 39200
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 6552 37120 6604 37126
rect 6552 37062 6604 37068
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 5724 36576 5776 36582
rect 5724 36518 5776 36524
rect 5736 32910 5764 36518
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 5828 32434 5856 37062
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 6564 31890 6592 37062
rect 6828 36032 6880 36038
rect 6828 35974 6880 35980
rect 6644 32768 6696 32774
rect 6644 32710 6696 32716
rect 6552 31884 6604 31890
rect 6552 31826 6604 31832
rect 5908 29164 5960 29170
rect 5908 29106 5960 29112
rect 5920 27130 5948 29106
rect 6000 27532 6052 27538
rect 6000 27474 6052 27480
rect 5908 27124 5960 27130
rect 5908 27066 5960 27072
rect 5816 26988 5868 26994
rect 6012 26976 6040 27474
rect 5816 26930 5868 26936
rect 5920 26948 6040 26976
rect 6460 26988 6512 26994
rect 5632 24880 5684 24886
rect 5632 24822 5684 24828
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5354 23080 5410 23089
rect 5354 23015 5410 23024
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 21944 5488 22918
rect 5552 22642 5580 24754
rect 5644 24206 5672 24822
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5644 23730 5672 24142
rect 5632 23724 5684 23730
rect 5684 23684 5764 23712
rect 5632 23666 5684 23672
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5460 21916 5580 21944
rect 5354 21720 5410 21729
rect 5354 21655 5410 21664
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5170 18864 5226 18873
rect 5170 18799 5226 18808
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 4908 17326 5028 17354
rect 4896 17128 4948 17134
rect 4894 17096 4896 17105
rect 4948 17096 4950 17105
rect 4894 17031 4950 17040
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4908 14414 4936 16662
rect 5000 15094 5028 17326
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16590 5120 16934
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4620 11824 4672 11830
rect 4526 11792 4582 11801
rect 4620 11766 4672 11772
rect 4526 11727 4582 11736
rect 4540 11694 4568 11727
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11218 4660 11766
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4264 10674 4292 11154
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9110 4660 11018
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 9104 4672 9110
rect 4066 9072 4122 9081
rect 4620 9046 4672 9052
rect 4724 9042 4752 9318
rect 4066 9007 4122 9016
rect 4712 9036 4764 9042
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3988 7970 4016 8434
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3896 7942 4016 7970
rect 3896 6866 3924 7942
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3528 2746 3648 2774
rect 3146 2680 3202 2689
rect 3146 2615 3202 2624
rect 3160 2446 3188 2615
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 1766 2136 1822 2145
rect 1766 2071 1822 2080
rect 1964 800 1992 2246
rect 3252 800 3280 2246
rect 3620 2038 3648 2746
rect 3608 2032 3660 2038
rect 3608 1974 3660 1980
rect 3712 1601 3740 4490
rect 3896 2553 3924 5238
rect 3988 3380 4016 7822
rect 4080 7342 4108 9007
rect 4712 8978 4764 8984
rect 4908 8974 4936 14350
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4540 7410 4568 7958
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6866 4660 8842
rect 5000 8820 5028 12582
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4908 8792 5028 8820
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4632 6225 4660 6666
rect 4618 6216 4674 6225
rect 4618 6151 4674 6160
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4436 5296 4488 5302
rect 4434 5264 4436 5273
rect 4488 5264 4490 5273
rect 4434 5199 4490 5208
rect 4540 5030 4568 5578
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4540 4049 4568 4762
rect 4526 4040 4582 4049
rect 4526 3975 4582 3984
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4080 3505 4108 3674
rect 4344 3664 4396 3670
rect 4342 3632 4344 3641
rect 4396 3632 4398 3641
rect 4342 3567 4398 3576
rect 4344 3528 4396 3534
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 4342 3496 4344 3505
rect 4396 3496 4398 3505
rect 4342 3431 4398 3440
rect 4436 3392 4488 3398
rect 3988 3352 4108 3380
rect 3882 2544 3938 2553
rect 3882 2479 3938 2488
rect 3884 2440 3936 2446
rect 4080 2417 4108 3352
rect 4632 3380 4660 5238
rect 4724 4758 4752 8502
rect 4802 7576 4858 7585
rect 4802 7511 4804 7520
rect 4856 7511 4858 7520
rect 4804 7482 4856 7488
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4321 4752 4558
rect 4710 4312 4766 4321
rect 4710 4247 4766 4256
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4488 3352 4660 3380
rect 4436 3334 4488 3340
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4448 2922 4476 3130
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4724 2774 4752 4014
rect 4816 3466 4844 7142
rect 4908 6118 4936 8792
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 5000 7954 5028 8366
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5000 7206 5028 7686
rect 5092 7342 5120 9862
rect 5184 9382 5212 18799
rect 5276 13954 5304 19178
rect 5368 15502 5396 21655
rect 5446 21312 5502 21321
rect 5446 21247 5502 21256
rect 5460 18290 5488 21247
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5448 17808 5500 17814
rect 5446 17776 5448 17785
rect 5500 17776 5502 17785
rect 5446 17711 5502 17720
rect 5446 17232 5502 17241
rect 5446 17167 5502 17176
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5460 14550 5488 17167
rect 5552 17082 5580 21916
rect 5644 17202 5672 23462
rect 5736 23118 5764 23684
rect 5828 23662 5856 26930
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5816 22976 5868 22982
rect 5816 22918 5868 22924
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5736 22545 5764 22578
rect 5722 22536 5778 22545
rect 5722 22471 5778 22480
rect 5722 21992 5778 22001
rect 5722 21927 5724 21936
rect 5776 21927 5778 21936
rect 5724 21898 5776 21904
rect 5722 21856 5778 21865
rect 5722 21791 5778 21800
rect 5736 19310 5764 21791
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18222 5764 19246
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5722 18048 5778 18057
rect 5722 17983 5778 17992
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5552 17054 5672 17082
rect 5644 16522 5672 17054
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5552 15638 5580 15982
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5736 14958 5764 17983
rect 5828 16182 5856 22918
rect 5920 22273 5948 26948
rect 6460 26930 6512 26936
rect 6472 26382 6500 26930
rect 6460 26376 6512 26382
rect 6458 26344 6460 26353
rect 6512 26344 6514 26353
rect 6458 26279 6514 26288
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6184 24744 6236 24750
rect 6184 24686 6236 24692
rect 6196 24410 6224 24686
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6000 23588 6052 23594
rect 6000 23530 6052 23536
rect 6012 22817 6040 23530
rect 6104 23497 6132 24142
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6184 23656 6236 23662
rect 6184 23598 6236 23604
rect 6090 23488 6146 23497
rect 6090 23423 6146 23432
rect 5998 22808 6054 22817
rect 5998 22743 6054 22752
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5906 22264 5962 22273
rect 5906 22199 5962 22208
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5920 20874 5948 21830
rect 6012 20874 6040 22578
rect 6092 22568 6144 22574
rect 6092 22510 6144 22516
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 5920 20398 5948 20810
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 5908 20392 5960 20398
rect 6012 20369 6040 20402
rect 5908 20334 5960 20340
rect 5998 20360 6054 20369
rect 5998 20295 6054 20304
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5276 13926 5396 13954
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 11642 5304 13806
rect 5368 13530 5396 13926
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5460 13326 5488 14350
rect 5644 14278 5672 14758
rect 5736 14482 5764 14894
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5920 13433 5948 17478
rect 6012 17377 6040 18566
rect 6104 18222 6132 22510
rect 6196 22438 6224 23598
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6182 22264 6238 22273
rect 6182 22199 6238 22208
rect 6196 21162 6224 22199
rect 6288 22137 6316 22578
rect 6274 22128 6330 22137
rect 6274 22063 6330 22072
rect 6274 21992 6330 22001
rect 6274 21927 6330 21936
rect 6288 21350 6316 21927
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6196 21134 6316 21162
rect 6182 21040 6238 21049
rect 6182 20975 6184 20984
rect 6236 20975 6238 20984
rect 6184 20946 6236 20952
rect 6184 20324 6236 20330
rect 6184 20266 6236 20272
rect 6196 19922 6224 20266
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6182 19816 6238 19825
rect 6182 19751 6184 19760
rect 6236 19751 6238 19760
rect 6184 19722 6236 19728
rect 6288 18601 6316 21134
rect 6274 18592 6330 18601
rect 6274 18527 6330 18536
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6104 17649 6132 18158
rect 6090 17640 6146 17649
rect 6090 17575 6146 17584
rect 5998 17368 6054 17377
rect 5998 17303 6054 17312
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6104 16794 6132 17274
rect 6380 16998 6408 23054
rect 6472 20369 6500 23666
rect 6564 23322 6592 24754
rect 6552 23316 6604 23322
rect 6552 23258 6604 23264
rect 6552 22024 6604 22030
rect 6550 21992 6552 22001
rect 6604 21992 6606 22001
rect 6550 21927 6606 21936
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 20806 6592 21830
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6458 20360 6514 20369
rect 6458 20295 6514 20304
rect 6564 19854 6592 20742
rect 6656 20534 6684 32710
rect 6736 31816 6788 31822
rect 6736 31758 6788 31764
rect 6748 29850 6776 31758
rect 6736 29844 6788 29850
rect 6736 29786 6788 29792
rect 6840 29170 6868 35974
rect 7852 32026 7880 37198
rect 9048 36922 9076 39200
rect 9404 37188 9456 37194
rect 9404 37130 9456 37136
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 9140 36378 9168 36722
rect 9128 36372 9180 36378
rect 9128 36314 9180 36320
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 9128 32224 9180 32230
rect 9128 32166 9180 32172
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 9036 31952 9088 31958
rect 9036 31894 9088 31900
rect 7656 31816 7708 31822
rect 7656 31758 7708 31764
rect 7668 31482 7696 31758
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7392 30433 7420 31282
rect 8576 30592 8628 30598
rect 8576 30534 8628 30540
rect 7378 30424 7434 30433
rect 7378 30359 7434 30368
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6828 29028 6880 29034
rect 6828 28970 6880 28976
rect 6736 26852 6788 26858
rect 6736 26794 6788 26800
rect 6748 25770 6776 26794
rect 6736 25764 6788 25770
rect 6736 25706 6788 25712
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6748 24886 6776 25094
rect 6736 24880 6788 24886
rect 6736 24822 6788 24828
rect 6840 23644 6868 28970
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7196 25832 7248 25838
rect 7196 25774 7248 25780
rect 7024 23730 7052 25774
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 6748 23616 6868 23644
rect 7024 23633 7052 23666
rect 7010 23624 7066 23633
rect 6748 20913 6776 23616
rect 7010 23559 7066 23568
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 6840 22642 6868 23054
rect 6920 23044 6972 23050
rect 6920 22986 6972 22992
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6932 22522 6960 22986
rect 6840 22494 6960 22522
rect 6840 21554 6868 22494
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6840 21457 6868 21490
rect 6826 21448 6882 21457
rect 6826 21383 6882 21392
rect 6734 20904 6790 20913
rect 6734 20839 6790 20848
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6458 17368 6514 17377
rect 6458 17303 6514 17312
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5538 13424 5594 13433
rect 5538 13359 5594 13368
rect 5906 13424 5962 13433
rect 5906 13359 5962 13368
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5552 12782 5580 13359
rect 5722 13288 5778 13297
rect 6012 13258 6040 16186
rect 6104 16130 6132 16730
rect 6104 16102 6316 16130
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6104 15638 6132 15846
rect 6092 15632 6144 15638
rect 6092 15574 6144 15580
rect 6196 15366 6224 15982
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6288 13870 6316 16102
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5722 13223 5778 13232
rect 6000 13252 6052 13258
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5448 12436 5500 12442
rect 5736 12434 5764 13223
rect 6000 13194 6052 13200
rect 6104 12986 6132 13466
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5448 12378 5500 12384
rect 5644 12406 5764 12434
rect 5356 12232 5408 12238
rect 5354 12200 5356 12209
rect 5408 12200 5410 12209
rect 5460 12186 5488 12378
rect 5460 12170 5580 12186
rect 5460 12164 5592 12170
rect 5460 12158 5540 12164
rect 5354 12135 5410 12144
rect 5540 12106 5592 12112
rect 5276 11614 5396 11642
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5276 11218 5304 11494
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5368 10554 5396 11614
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5276 10526 5396 10554
rect 5276 10470 5304 10526
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5276 7546 5304 9862
rect 5446 9752 5502 9761
rect 5446 9687 5502 9696
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 5000 5778 5028 6666
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4896 4684 4948 4690
rect 5000 4672 5028 5714
rect 5276 5250 5304 7346
rect 4948 4644 5028 4672
rect 5092 5222 5304 5250
rect 4896 4626 4948 4632
rect 4908 4282 4936 4626
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5092 4434 5120 5222
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5184 4554 5212 5102
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5276 4486 5304 4966
rect 5368 4826 5396 7482
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5460 4706 5488 9687
rect 5552 9518 5580 11494
rect 5644 10266 5672 12406
rect 5906 11928 5962 11937
rect 5906 11863 5962 11872
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5552 8566 5580 9454
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5552 7410 5580 8366
rect 5644 8022 5672 8842
rect 5736 8430 5764 11290
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5736 7886 5764 8230
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5828 7546 5856 11154
rect 5920 10130 5948 11863
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5920 9722 5948 9930
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5920 9110 5948 9522
rect 6012 9518 6040 12786
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5920 7886 5948 8910
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5920 7478 5948 7822
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5368 4678 5488 4706
rect 5264 4480 5316 4486
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4908 3398 4936 4218
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2746 4752 2774
rect 3884 2382 3936 2388
rect 4066 2408 4122 2417
rect 3698 1592 3754 1601
rect 3698 1527 3754 1536
rect 3896 800 3924 2382
rect 4632 2378 4660 2746
rect 4066 2343 4122 2352
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 5000 1222 5028 4422
rect 5092 4406 5212 4434
rect 5264 4422 5316 4428
rect 5078 4312 5134 4321
rect 5078 4247 5080 4256
rect 5132 4247 5134 4256
rect 5080 4218 5132 4224
rect 5078 4040 5134 4049
rect 5078 3975 5134 3984
rect 5092 3097 5120 3975
rect 5078 3088 5134 3097
rect 5184 3058 5212 4406
rect 5276 4078 5304 4422
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5078 3023 5134 3032
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5184 2961 5212 2994
rect 5170 2952 5226 2961
rect 5170 2887 5226 2896
rect 5368 2774 5396 4678
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5460 3194 5488 4490
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5552 3126 5580 5646
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5644 2990 5672 5782
rect 5722 5128 5778 5137
rect 5722 5063 5724 5072
rect 5776 5063 5778 5072
rect 5724 5034 5776 5040
rect 5722 4584 5778 4593
rect 5722 4519 5778 4528
rect 5736 4146 5764 4519
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5736 2854 5764 4082
rect 5828 3233 5856 7346
rect 5920 6798 5948 7414
rect 6012 7002 6040 9454
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 6458 5948 6734
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 4078 6040 6054
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6104 3738 6132 9862
rect 6182 6896 6238 6905
rect 6182 6831 6238 6840
rect 6196 4146 6224 6831
rect 6380 6474 6408 16730
rect 6472 15434 6500 17303
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 14006 6500 14418
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6564 13394 6592 18702
rect 6656 14362 6684 20266
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6748 18358 6776 20198
rect 6840 18873 6868 21383
rect 6932 20482 6960 22374
rect 7012 21956 7064 21962
rect 7012 21898 7064 21904
rect 7024 20777 7052 21898
rect 7010 20768 7066 20777
rect 7010 20703 7066 20712
rect 7116 20534 7144 24006
rect 7208 21622 7236 25774
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7196 21616 7248 21622
rect 7300 21604 7328 22374
rect 7484 22137 7512 22918
rect 7470 22128 7526 22137
rect 7470 22063 7526 22072
rect 7576 21978 7604 24550
rect 7852 24410 7880 26862
rect 8024 26784 8076 26790
rect 8024 26726 8076 26732
rect 8036 25906 8064 26726
rect 8024 25900 8076 25906
rect 8024 25842 8076 25848
rect 7932 25832 7984 25838
rect 7932 25774 7984 25780
rect 7944 25362 7972 25774
rect 7932 25356 7984 25362
rect 7932 25298 7984 25304
rect 8116 24880 8168 24886
rect 8116 24822 8168 24828
rect 7932 24676 7984 24682
rect 7932 24618 7984 24624
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7852 23730 7880 24346
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7484 21950 7604 21978
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7380 21616 7432 21622
rect 7300 21576 7380 21604
rect 7196 21558 7248 21564
rect 7380 21558 7432 21564
rect 7288 21412 7340 21418
rect 7288 21354 7340 21360
rect 7300 21026 7328 21354
rect 7484 21078 7512 21950
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7208 20998 7328 21026
rect 7472 21072 7524 21078
rect 7472 21014 7524 21020
rect 7104 20528 7156 20534
rect 6932 20454 7052 20482
rect 7104 20470 7156 20476
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 19990 6960 20334
rect 7024 20262 7052 20454
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 7024 19417 7052 19722
rect 7010 19408 7066 19417
rect 7010 19343 7066 19352
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6826 18864 6882 18873
rect 6826 18799 6882 18808
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6840 18426 6868 18702
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6932 18222 6960 19246
rect 7102 19136 7158 19145
rect 7102 19071 7158 19080
rect 7116 18698 7144 19071
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7116 18601 7144 18634
rect 7102 18592 7158 18601
rect 7102 18527 7158 18536
rect 7010 18320 7066 18329
rect 7010 18255 7066 18264
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6932 18034 6960 18158
rect 6840 18006 6960 18034
rect 6840 17746 6868 18006
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6734 17096 6790 17105
rect 6734 17031 6790 17040
rect 6748 16998 6776 17031
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6840 15570 6868 17682
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6748 14498 6776 15370
rect 6840 14958 6868 15506
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6748 14470 6868 14498
rect 6656 14346 6776 14362
rect 6656 14340 6788 14346
rect 6656 14334 6736 14340
rect 6736 14282 6788 14288
rect 6840 13954 6868 14470
rect 6656 13926 6868 13954
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6656 12434 6684 13926
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6472 12406 6684 12434
rect 6472 10962 6500 12406
rect 6748 12322 6776 13738
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 12617 6868 12854
rect 6826 12608 6882 12617
rect 6826 12543 6882 12552
rect 6656 12294 6776 12322
rect 6472 10934 6592 10962
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6472 9042 6500 10746
rect 6564 9586 6592 10934
rect 6656 10810 6684 12294
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6748 11830 6776 12174
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6932 11370 6960 15302
rect 7024 14890 7052 18255
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7116 16658 7144 17070
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 16114 7144 16594
rect 7208 16561 7236 20998
rect 7576 20874 7604 21830
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7300 19446 7328 20810
rect 7668 19786 7696 21966
rect 7852 21944 7880 23530
rect 7944 23322 7972 24618
rect 8022 24168 8078 24177
rect 8022 24103 8078 24112
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7760 21916 7880 21944
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7470 19544 7526 19553
rect 7470 19479 7526 19488
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 7286 19000 7342 19009
rect 7286 18935 7342 18944
rect 7194 16552 7250 16561
rect 7194 16487 7250 16496
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7102 15056 7158 15065
rect 7102 14991 7104 15000
rect 7156 14991 7158 15000
rect 7104 14962 7156 14968
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7208 14618 7236 15642
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13938 7236 14214
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 13326 7236 13670
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12850 7144 13126
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7010 12472 7066 12481
rect 7010 12407 7066 12416
rect 7024 12306 7052 12407
rect 7116 12306 7144 12786
rect 7300 12646 7328 18935
rect 7380 18692 7432 18698
rect 7380 18634 7432 18640
rect 7392 14006 7420 18634
rect 7484 18630 7512 19479
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7484 15026 7512 18566
rect 7654 16552 7710 16561
rect 7654 16487 7656 16496
rect 7708 16487 7710 16496
rect 7656 16458 7708 16464
rect 7654 16280 7710 16289
rect 7654 16215 7710 16224
rect 7668 16182 7696 16215
rect 7656 16176 7708 16182
rect 7656 16118 7708 16124
rect 7760 15366 7788 21916
rect 7838 21856 7894 21865
rect 7838 21791 7894 21800
rect 7852 15434 7880 21791
rect 7944 20602 7972 23258
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 8036 19174 8064 24103
rect 8128 22778 8156 24822
rect 8220 24750 8248 27066
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8312 24206 8340 25638
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 8036 16454 8064 19110
rect 8128 18737 8156 21966
rect 8114 18728 8170 18737
rect 8114 18663 8170 18672
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 8128 16266 8156 18663
rect 8036 16238 8156 16266
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 8036 15178 8064 16238
rect 8114 15600 8170 15609
rect 8114 15535 8170 15544
rect 7760 15150 8064 15178
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7484 14906 7512 14962
rect 7484 14878 7604 14906
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 14006 7512 14758
rect 7576 14414 7604 14878
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7484 12434 7512 13806
rect 7300 12406 7512 12434
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6748 11354 6960 11370
rect 6736 11348 6960 11354
rect 6788 11342 6960 11348
rect 6736 11290 6788 11296
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6828 10736 6880 10742
rect 6826 10704 6828 10713
rect 6880 10704 6882 10713
rect 6826 10639 6882 10648
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6656 10266 6684 10406
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6828 10124 6880 10130
rect 6880 10084 6960 10112
rect 6828 10066 6880 10072
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6550 9480 6606 9489
rect 6550 9415 6552 9424
rect 6604 9415 6606 9424
rect 6552 9386 6604 9392
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6564 8294 6592 8978
rect 6656 8786 6684 9998
rect 6932 9518 6960 10084
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6734 8936 6790 8945
rect 6734 8871 6736 8880
rect 6788 8871 6790 8880
rect 6736 8842 6788 8848
rect 6656 8758 6776 8786
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 7834 6684 7890
rect 6472 7818 6684 7834
rect 6460 7812 6684 7818
rect 6512 7806 6684 7812
rect 6460 7754 6512 7760
rect 6288 6446 6408 6474
rect 6288 5166 6316 6446
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5814 3224 5870 3233
rect 5814 3159 5870 3168
rect 5828 3058 5856 3159
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6380 2854 6408 6326
rect 6472 5914 6500 7754
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6564 7313 6592 7346
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6564 6866 6592 7239
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6564 5234 6592 6122
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6472 2990 6500 4150
rect 6564 3505 6592 5170
rect 6656 5166 6684 7346
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6748 4049 6776 8758
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 6882 6960 7278
rect 6840 6854 6960 6882
rect 6840 6322 6868 6854
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 5710 6868 6258
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5370 6868 5646
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6840 4214 6868 5306
rect 6918 5264 6974 5273
rect 6918 5199 6974 5208
rect 6932 4486 6960 5199
rect 7024 4622 7052 11698
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6734 4040 6790 4049
rect 6644 4004 6696 4010
rect 6734 3975 6790 3984
rect 6644 3946 6696 3952
rect 6550 3496 6606 3505
rect 6656 3466 6684 3946
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3602 6776 3878
rect 6826 3632 6882 3641
rect 6736 3596 6788 3602
rect 6826 3567 6882 3576
rect 6736 3538 6788 3544
rect 6840 3534 6868 3567
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6550 3431 6606 3440
rect 6644 3460 6696 3466
rect 6564 3058 6592 3431
rect 6644 3402 6696 3408
rect 6644 3120 6696 3126
rect 6932 3108 6960 4150
rect 7024 3670 7052 4558
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6696 3080 6960 3108
rect 6644 3062 6696 3068
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 5368 2746 5488 2774
rect 5460 2582 5488 2746
rect 7024 2650 7052 3334
rect 7116 2774 7144 10406
rect 7208 7002 7236 11018
rect 7300 10674 7328 12406
rect 7484 12345 7512 12406
rect 7470 12336 7526 12345
rect 7470 12271 7526 12280
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7562 11384 7618 11393
rect 7668 11354 7696 11562
rect 7562 11319 7564 11328
rect 7616 11319 7618 11328
rect 7656 11348 7708 11354
rect 7564 11290 7616 11296
rect 7656 11290 7708 11296
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 10470 7328 10610
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7392 8514 7420 11018
rect 7760 10826 7788 15150
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7852 14618 7880 15030
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8036 14414 8064 14554
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 12646 7880 13806
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 11830 7880 12582
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7576 10798 7788 10826
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 10130 7512 10406
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7300 8486 7420 8514
rect 7300 8106 7328 8486
rect 7484 8430 7512 9454
rect 7576 9110 7604 10798
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7760 10130 7788 10678
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7852 10169 7880 10474
rect 7838 10160 7894 10169
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7748 10124 7800 10130
rect 7838 10095 7894 10104
rect 7748 10066 7800 10072
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7392 8242 7420 8298
rect 7576 8242 7604 9046
rect 7392 8214 7604 8242
rect 7300 8078 7420 8106
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7194 6488 7250 6497
rect 7194 6423 7250 6432
rect 7208 6390 7236 6423
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7208 6089 7236 6326
rect 7194 6080 7250 6089
rect 7194 6015 7250 6024
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 5642 7236 5714
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7392 4185 7420 8078
rect 7668 8022 7696 10066
rect 7944 9976 7972 12854
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 11286 8064 12242
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 8036 10742 8064 11222
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7760 9948 7972 9976
rect 7760 9178 7788 9948
rect 8128 9874 8156 15535
rect 8220 13258 8248 22918
rect 8298 22536 8354 22545
rect 8298 22471 8354 22480
rect 8312 21894 8340 22471
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8404 20942 8432 22102
rect 8392 20936 8444 20942
rect 8298 20904 8354 20913
rect 8392 20878 8444 20884
rect 8298 20839 8300 20848
rect 8352 20839 8354 20848
rect 8300 20810 8352 20816
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 13297 8340 20198
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8404 19553 8432 19858
rect 8390 19544 8446 19553
rect 8390 19479 8446 19488
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 15337 8432 19110
rect 8496 15366 8524 25230
rect 8588 23798 8616 30534
rect 8944 29640 8996 29646
rect 8944 29582 8996 29588
rect 8956 27062 8984 29582
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8956 24682 8984 26998
rect 8944 24676 8996 24682
rect 8944 24618 8996 24624
rect 8576 23792 8628 23798
rect 8576 23734 8628 23740
rect 8668 23588 8720 23594
rect 8668 23530 8720 23536
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8588 22642 8616 23054
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8588 18970 8616 22578
rect 8680 21010 8708 23530
rect 8852 23248 8904 23254
rect 8852 23190 8904 23196
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8668 21004 8720 21010
rect 8668 20946 8720 20952
rect 8772 20534 8800 22374
rect 8864 21486 8892 23190
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8864 20602 8892 21422
rect 8956 21146 8984 21422
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 8956 19718 8984 21082
rect 9048 20398 9076 31894
rect 9140 24138 9168 32166
rect 9324 27452 9352 32302
rect 9416 30734 9444 37130
rect 9692 37126 9720 39200
rect 10980 37330 11008 39200
rect 10968 37324 11020 37330
rect 10968 37266 11020 37272
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 11796 37256 11848 37262
rect 12268 37244 12296 39200
rect 12440 37256 12492 37262
rect 12268 37216 12440 37244
rect 11796 37198 11848 37204
rect 12440 37198 12492 37204
rect 9680 37120 9732 37126
rect 9680 37062 9732 37068
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9784 30297 9812 37198
rect 11808 31754 11836 37198
rect 13556 37126 13584 39200
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 11624 31726 11836 31754
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 9770 30288 9826 30297
rect 9770 30223 9826 30232
rect 10600 29504 10652 29510
rect 10600 29446 10652 29452
rect 9324 27424 9444 27452
rect 9312 26512 9364 26518
rect 9312 26454 9364 26460
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 9232 25294 9260 25978
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9324 24886 9352 26454
rect 9416 25906 9444 27424
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9588 26308 9640 26314
rect 9588 26250 9640 26256
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9312 24880 9364 24886
rect 9312 24822 9364 24828
rect 9416 24750 9444 25842
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 9232 24274 9260 24686
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9128 24132 9180 24138
rect 9128 24074 9180 24080
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9140 20262 9168 22578
rect 9218 22536 9274 22545
rect 9218 22471 9274 22480
rect 9232 21962 9260 22471
rect 9324 21962 9352 22918
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9312 21956 9364 21962
rect 9312 21898 9364 21904
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9324 21146 9352 21354
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8588 17134 8616 18906
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8484 15360 8536 15366
rect 8390 15328 8446 15337
rect 8484 15302 8536 15308
rect 8390 15263 8446 15272
rect 8496 15162 8524 15302
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 13326 8432 14214
rect 8392 13320 8444 13326
rect 8298 13288 8354 13297
rect 8208 13252 8260 13258
rect 8392 13262 8444 13268
rect 8298 13223 8354 13232
rect 8208 13194 8260 13200
rect 8404 11218 8432 13262
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 11830 8524 13126
rect 8588 12481 8616 16526
rect 8680 14550 8708 18906
rect 8944 18896 8996 18902
rect 8850 18864 8906 18873
rect 8944 18838 8996 18844
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 8850 18799 8906 18808
rect 8864 18204 8892 18799
rect 8956 18601 8984 18838
rect 8942 18592 8998 18601
rect 8942 18527 8998 18536
rect 8944 18216 8996 18222
rect 8864 18176 8944 18204
rect 8758 15464 8814 15473
rect 8758 15399 8814 15408
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8574 12472 8630 12481
rect 8574 12407 8630 12416
rect 8588 12238 8616 12407
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8680 11354 8708 12718
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7852 9846 8156 9874
rect 7852 9518 7880 9846
rect 8220 9674 8248 11086
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8404 10198 8432 10678
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8482 10160 8538 10169
rect 8482 10095 8538 10104
rect 8496 9926 8524 10095
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8024 9648 8076 9654
rect 8220 9646 8340 9674
rect 8076 9608 8156 9636
rect 8024 9590 8076 9596
rect 8128 9518 8156 9608
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7760 8634 7788 8842
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7654 7168 7710 7177
rect 7654 7103 7710 7112
rect 7668 7002 7696 7103
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7576 6662 7604 6938
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7378 4176 7434 4185
rect 7378 4111 7434 4120
rect 7576 3194 7604 5578
rect 7852 5166 7880 9318
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7746 4992 7802 5001
rect 7746 4927 7802 4936
rect 7760 4622 7788 4927
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7668 3534 7696 4014
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7852 3233 7880 4558
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7838 3224 7894 3233
rect 7564 3188 7616 3194
rect 7838 3159 7894 3168
rect 7564 3130 7616 3136
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7208 2922 7236 3062
rect 7852 3058 7880 3159
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7392 2961 7420 2994
rect 7944 2990 7972 4422
rect 8036 3233 8064 8910
rect 8312 8072 8340 9646
rect 8772 8838 8800 15399
rect 8864 14521 8892 18176
rect 8944 18158 8996 18164
rect 8942 17776 8998 17785
rect 8942 17711 8944 17720
rect 8996 17711 8998 17720
rect 8944 17682 8996 17688
rect 8850 14512 8906 14521
rect 8850 14447 8906 14456
rect 8864 14414 8892 14447
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8850 13832 8906 13841
rect 8850 13767 8906 13776
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8128 8044 8340 8072
rect 8128 7410 8156 8044
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8220 7002 8248 7754
rect 8312 7206 8340 7890
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7546 8432 7686
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8128 5846 8156 6666
rect 8220 6254 8248 6734
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8404 5574 8432 5850
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8022 3224 8078 3233
rect 8128 3194 8156 5510
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8404 4622 8432 4762
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8312 3534 8340 4082
rect 8496 3738 8524 8502
rect 8574 8256 8630 8265
rect 8574 8191 8630 8200
rect 8588 7478 8616 8191
rect 8864 7954 8892 13767
rect 9048 13462 9076 18838
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 16697 9168 17478
rect 9126 16688 9182 16697
rect 9126 16623 9182 16632
rect 9232 15994 9260 20810
rect 9416 19786 9444 22374
rect 9508 21350 9536 23122
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9600 21146 9628 26250
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9692 23866 9720 25094
rect 9784 24070 9812 27338
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 10060 26450 10088 26726
rect 10140 26512 10192 26518
rect 10140 26454 10192 26460
rect 10048 26444 10100 26450
rect 10048 26386 10100 26392
rect 10152 25702 10180 26454
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 10232 25696 10284 25702
rect 10232 25638 10284 25644
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9784 23730 9812 24006
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9692 20806 9720 22986
rect 9784 21622 9812 23462
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 10060 22778 10088 22986
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 9968 22438 9996 22714
rect 10152 22710 10180 25094
rect 10244 24138 10272 25638
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10232 24132 10284 24138
rect 10232 24074 10284 24080
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 10232 22704 10284 22710
rect 10232 22646 10284 22652
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9876 22234 9904 22374
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9784 20482 9812 20946
rect 9876 20874 9904 21558
rect 9954 21312 10010 21321
rect 9954 21247 10010 21256
rect 9968 21078 9996 21247
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9692 20454 9812 20482
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9508 19990 9536 20266
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9324 18358 9352 19110
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9324 17066 9352 17546
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 9416 16969 9444 18566
rect 9402 16960 9458 16969
rect 9402 16895 9458 16904
rect 9600 16833 9628 18634
rect 9692 17320 9720 20454
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9784 19922 9812 20334
rect 9862 19952 9918 19961
rect 9772 19916 9824 19922
rect 9862 19887 9918 19896
rect 9772 19858 9824 19864
rect 9876 19334 9904 19887
rect 9956 19440 10008 19446
rect 9954 19408 9956 19417
rect 10008 19408 10010 19417
rect 9954 19343 10010 19352
rect 9784 19306 9904 19334
rect 9784 17785 9812 19306
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9862 18456 9918 18465
rect 9862 18391 9918 18400
rect 9876 18222 9904 18391
rect 9968 18222 9996 18906
rect 10060 18766 10088 22034
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 18358 10088 18566
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9770 17776 9826 17785
rect 9770 17711 9826 17720
rect 10048 17332 10100 17338
rect 9692 17292 9904 17320
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9310 16824 9366 16833
rect 9310 16759 9312 16768
rect 9364 16759 9366 16768
rect 9586 16824 9642 16833
rect 9586 16759 9642 16768
rect 9312 16730 9364 16736
rect 9588 16720 9640 16726
rect 9310 16688 9366 16697
rect 9416 16680 9588 16708
rect 9416 16674 9444 16680
rect 9366 16646 9444 16674
rect 9588 16662 9640 16668
rect 9310 16623 9366 16632
rect 9140 15966 9260 15994
rect 9140 15910 9168 15966
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9126 15328 9182 15337
rect 9126 15263 9182 15272
rect 9140 15162 9168 15263
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 8956 12714 8984 13330
rect 9048 13258 9076 13398
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9140 12850 9168 13330
rect 9232 12918 9260 15846
rect 9324 15201 9352 16623
rect 9588 16584 9640 16590
rect 9586 16552 9588 16561
rect 9640 16552 9642 16561
rect 9692 16522 9720 17138
rect 9586 16487 9642 16496
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 16250 9628 16390
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9310 15192 9366 15201
rect 9310 15127 9366 15136
rect 9494 14376 9550 14385
rect 9404 14340 9456 14346
rect 9494 14311 9496 14320
rect 9404 14282 9456 14288
rect 9548 14311 9550 14320
rect 9496 14282 9548 14288
rect 9416 13870 9444 14282
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9508 13530 9536 13874
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9404 13388 9456 13394
rect 9324 13348 9404 13376
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 9140 12646 9168 12786
rect 9324 12782 9352 13348
rect 9404 13330 9456 13336
rect 9600 13190 9628 15302
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9586 13016 9642 13025
rect 9586 12951 9642 12960
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9312 12436 9364 12442
rect 9508 12434 9536 12582
rect 9312 12378 9364 12384
rect 9416 12406 9536 12434
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9048 11898 9076 12106
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9324 11393 9352 12378
rect 9310 11384 9366 11393
rect 9310 11319 9366 11328
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 6905 8616 7278
rect 8574 6896 8630 6905
rect 8574 6831 8630 6840
rect 8574 6216 8630 6225
rect 8574 6151 8630 6160
rect 8588 5710 8616 6151
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8588 3670 8616 5170
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8022 3159 8078 3168
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 7932 2984 7984 2990
rect 7378 2952 7434 2961
rect 7196 2916 7248 2922
rect 7932 2926 7984 2932
rect 7378 2887 7434 2896
rect 7196 2858 7248 2864
rect 7116 2746 7236 2774
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 7208 2446 7236 2746
rect 8220 2446 8248 2994
rect 8312 2582 8340 3470
rect 8680 3398 8708 7686
rect 8850 7304 8906 7313
rect 8850 7239 8906 7248
rect 8758 7168 8814 7177
rect 8758 7103 8814 7112
rect 8772 6934 8800 7103
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8864 6866 8892 7239
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8956 5114 8984 11154
rect 9048 7834 9076 11154
rect 9232 8566 9260 11222
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9324 8430 9352 11319
rect 9416 8634 9444 12406
rect 9600 9738 9628 12951
rect 9692 12918 9720 16458
rect 9770 16144 9826 16153
rect 9770 16079 9772 16088
rect 9824 16079 9826 16088
rect 9772 16050 9824 16056
rect 9876 15978 9904 17292
rect 10048 17274 10100 17280
rect 10060 17202 10088 17274
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9968 15162 9996 16730
rect 10152 16590 10180 19722
rect 10244 19310 10272 22646
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10230 18864 10286 18873
rect 10230 18799 10286 18808
rect 10244 17513 10272 18799
rect 10230 17504 10286 17513
rect 10230 17439 10286 17448
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10244 16402 10272 17439
rect 10060 16374 10272 16402
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9784 12764 9812 14758
rect 9968 14618 9996 14894
rect 10060 14822 10088 16374
rect 10336 16130 10364 23666
rect 10520 22556 10548 24346
rect 10428 22528 10548 22556
rect 10428 19281 10456 22528
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10520 21593 10548 22374
rect 10612 22094 10640 29446
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11072 26994 11100 27270
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 10876 26920 10928 26926
rect 10876 26862 10928 26868
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10888 26518 10916 26862
rect 10876 26512 10928 26518
rect 10876 26454 10928 26460
rect 10980 26450 11008 26862
rect 10968 26444 11020 26450
rect 10968 26386 11020 26392
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 11164 26246 11192 26318
rect 11152 26240 11204 26246
rect 11152 26182 11204 26188
rect 11256 26024 11284 27814
rect 11164 25996 11284 26024
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10796 25430 10824 25842
rect 10784 25424 10836 25430
rect 10784 25366 10836 25372
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10704 22710 10732 24074
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10796 22574 10824 25162
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10980 24206 11008 24754
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10784 22568 10836 22574
rect 10782 22536 10784 22545
rect 10836 22536 10838 22545
rect 10782 22471 10838 22480
rect 10612 22066 10732 22094
rect 10506 21584 10562 21593
rect 10506 21519 10562 21528
rect 10600 21548 10652 21554
rect 10520 20534 10548 21519
rect 10600 21490 10652 21496
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10612 19334 10640 21490
rect 10520 19306 10640 19334
rect 10414 19272 10470 19281
rect 10414 19207 10470 19216
rect 10520 18850 10548 19306
rect 10428 18822 10548 18850
rect 10428 16289 10456 18822
rect 10508 18760 10560 18766
rect 10560 18720 10640 18748
rect 10508 18702 10560 18708
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10520 16425 10548 16526
rect 10506 16416 10562 16425
rect 10506 16351 10562 16360
rect 10414 16280 10470 16289
rect 10414 16215 10470 16224
rect 10244 16102 10364 16130
rect 10520 16114 10548 16351
rect 10416 16108 10468 16114
rect 10244 15094 10272 16102
rect 10416 16050 10468 16056
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15910 10364 15982
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15434 10364 15846
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9692 12736 9812 12764
rect 9692 11665 9720 12736
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9678 11656 9734 11665
rect 9678 11591 9734 11600
rect 9692 11558 9720 11591
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10470 9720 11086
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9784 9926 9812 12106
rect 9876 11762 9904 14554
rect 9968 13530 9996 14554
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 10060 14006 10088 14039
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 10060 13870 10088 13942
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9968 11898 9996 12650
rect 10060 12170 10088 12854
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9954 11520 10010 11529
rect 9954 11455 10010 11464
rect 9968 11354 9996 11455
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 10152 10674 10180 14826
rect 10244 13802 10272 15030
rect 10428 14550 10456 16050
rect 10520 14890 10548 16050
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10428 14362 10456 14486
rect 10428 14334 10548 14362
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 10244 12345 10272 12951
rect 10230 12336 10286 12345
rect 10230 12271 10286 12280
rect 10244 12238 10272 12271
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10336 11354 10364 14214
rect 10428 14006 10456 14214
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10520 13938 10548 14334
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10612 13025 10640 18720
rect 10704 18698 10732 22066
rect 10782 21992 10838 22001
rect 10888 21962 10916 23462
rect 10782 21927 10784 21936
rect 10836 21927 10838 21936
rect 10876 21956 10928 21962
rect 10784 21898 10836 21904
rect 10876 21898 10928 21904
rect 10796 21729 10824 21898
rect 10782 21720 10838 21729
rect 10782 21655 10838 21664
rect 10980 21434 11008 24142
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11072 21865 11100 23666
rect 11164 23186 11192 25996
rect 11348 25362 11376 30534
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 11058 21856 11114 21865
rect 11114 21814 11192 21842
rect 11058 21791 11114 21800
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10796 21406 11008 21434
rect 10796 19122 10824 21406
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10888 20534 10916 21286
rect 10966 21040 11022 21049
rect 10966 20975 10968 20984
rect 11020 20975 11022 20984
rect 10968 20946 11020 20952
rect 11072 20777 11100 21626
rect 11164 21486 11192 21814
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11058 20768 11114 20777
rect 11058 20703 11114 20712
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10888 20058 10916 20198
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10966 19680 11022 19689
rect 10966 19615 11022 19624
rect 10980 19514 11008 19615
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10796 19094 10916 19122
rect 10888 18873 10916 19094
rect 10874 18864 10930 18873
rect 10874 18799 10930 18808
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10704 18222 10732 18634
rect 10796 18290 10824 18634
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10876 18080 10928 18086
rect 10980 18068 11008 19178
rect 11072 19009 11100 19246
rect 11058 19000 11114 19009
rect 11058 18935 11114 18944
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 10928 18040 11008 18068
rect 10876 18022 10928 18028
rect 10704 17270 10732 18022
rect 10888 17921 10916 18022
rect 10874 17912 10930 17921
rect 10784 17876 10836 17882
rect 10874 17847 10930 17856
rect 10784 17818 10836 17824
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10704 15570 10732 17206
rect 10796 16250 10824 17818
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10876 17536 10928 17542
rect 10874 17504 10876 17513
rect 10928 17504 10930 17513
rect 10874 17439 10930 17448
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16969 10916 17070
rect 10874 16960 10930 16969
rect 10874 16895 10930 16904
rect 10980 16697 11008 17546
rect 11072 16726 11100 18294
rect 11060 16720 11112 16726
rect 10966 16688 11022 16697
rect 11060 16662 11112 16668
rect 10966 16623 11022 16632
rect 11164 16522 11192 20878
rect 11256 20602 11284 24006
rect 11348 21078 11376 25298
rect 11440 25226 11468 25638
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11440 21690 11468 21898
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11336 21072 11388 21078
rect 11336 21014 11388 21020
rect 11440 20641 11468 21626
rect 11532 21298 11560 22578
rect 11624 21622 11652 31726
rect 12360 30258 12388 37062
rect 14200 36854 14228 39200
rect 15488 37262 15516 39200
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 15476 37256 15528 37262
rect 15476 37198 15528 37204
rect 14292 36922 14320 37198
rect 15568 37120 15620 37126
rect 15568 37062 15620 37068
rect 14280 36916 14332 36922
rect 14280 36858 14332 36864
rect 14188 36848 14240 36854
rect 14188 36790 14240 36796
rect 13544 36780 13596 36786
rect 13544 36722 13596 36728
rect 15384 36780 15436 36786
rect 15384 36722 15436 36728
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 11992 26790 12020 27406
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11888 26512 11940 26518
rect 11888 26454 11940 26460
rect 11900 25498 11928 26454
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11704 24676 11756 24682
rect 11704 24618 11756 24624
rect 11612 21616 11664 21622
rect 11612 21558 11664 21564
rect 11532 21270 11652 21298
rect 11518 21176 11574 21185
rect 11518 21111 11520 21120
rect 11572 21111 11574 21120
rect 11520 21082 11572 21088
rect 11426 20632 11482 20641
rect 11244 20596 11296 20602
rect 11426 20567 11482 20576
rect 11244 20538 11296 20544
rect 11426 20088 11482 20097
rect 11426 20023 11482 20032
rect 11440 19378 11468 20023
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11532 19689 11560 19722
rect 11518 19680 11574 19689
rect 11518 19615 11574 19624
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11624 18986 11652 21270
rect 11348 18958 11652 18986
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14414 10824 14758
rect 10692 14408 10744 14414
rect 10690 14376 10692 14385
rect 10784 14408 10836 14414
rect 10744 14376 10746 14385
rect 10784 14350 10836 14356
rect 10690 14311 10746 14320
rect 10888 14260 10916 16390
rect 10966 15872 11022 15881
rect 10966 15807 11022 15816
rect 10704 14232 10916 14260
rect 10598 13016 10654 13025
rect 10598 12951 10654 12960
rect 10704 12442 10732 14232
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10414 12336 10470 12345
rect 10414 12271 10470 12280
rect 10428 11626 10456 12271
rect 10796 12050 10824 13874
rect 10520 12022 10824 12050
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 9680 9920 9732 9926
rect 9678 9888 9680 9897
rect 9772 9920 9824 9926
rect 9732 9888 9734 9897
rect 9772 9862 9824 9868
rect 9678 9823 9734 9832
rect 9508 9710 9628 9738
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9312 8424 9364 8430
rect 9218 8392 9274 8401
rect 9128 8356 9180 8362
rect 9312 8366 9364 8372
rect 9218 8327 9274 8336
rect 9128 8298 9180 8304
rect 9140 7954 9168 8298
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9048 7806 9168 7834
rect 9034 6896 9090 6905
rect 9034 6831 9090 6840
rect 9048 6798 9076 6831
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8864 5086 8984 5114
rect 8864 4146 8892 5086
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 4690 8984 4966
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8208 2440 8260 2446
rect 8484 2440 8536 2446
rect 8208 2382 8260 2388
rect 8404 2400 8484 2428
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 4988 1216 5040 1222
rect 4988 1158 5040 1164
rect 5184 800 5212 2246
rect 5276 1873 5304 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 5262 1864 5318 1873
rect 5262 1799 5318 1808
rect 6472 800 6500 2246
rect 6564 2009 6592 2382
rect 6550 2000 6606 2009
rect 6550 1935 6606 1944
rect 7116 870 7236 898
rect 7116 800 7144 870
rect 1398 776 1454 785
rect 1398 711 1454 720
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 7208 66 7236 870
rect 8404 800 8432 2400
rect 8484 2382 8536 2388
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8588 1834 8616 2314
rect 9048 1902 9076 6326
rect 9140 4078 9168 7806
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9232 2514 9260 8327
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9324 7818 9352 8230
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9416 7546 9444 7754
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9404 6792 9456 6798
rect 9402 6760 9404 6769
rect 9456 6760 9458 6769
rect 9402 6695 9458 6704
rect 9508 6610 9536 9710
rect 9588 9648 9640 9654
rect 9586 9616 9588 9625
rect 9640 9616 9642 9625
rect 9784 9586 9812 9862
rect 10244 9674 10272 10610
rect 10520 10470 10548 12022
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10612 10985 10640 11086
rect 10598 10976 10654 10985
rect 10598 10911 10654 10920
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10520 9722 10548 9862
rect 9876 9646 10272 9674
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 9586 9551 9642 9560
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9678 8256 9734 8265
rect 9678 8191 9734 8200
rect 9586 7032 9642 7041
rect 9586 6967 9642 6976
rect 9600 6662 9628 6967
rect 9692 6934 9720 8191
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9784 6866 9812 9522
rect 9876 8974 9904 9646
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 8974 10180 9318
rect 10428 9042 10456 9386
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9876 8514 9904 8910
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8634 9996 8774
rect 10414 8664 10470 8673
rect 9956 8628 10008 8634
rect 10414 8599 10470 8608
rect 9956 8570 10008 8576
rect 9876 8486 9996 8514
rect 10428 8498 10456 8599
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9416 6582 9536 6610
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9416 6390 9444 6582
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9324 6236 9352 6326
rect 9692 6236 9720 6734
rect 9324 6208 9720 6236
rect 9692 5030 9720 6208
rect 9784 5642 9812 6802
rect 9876 6390 9904 7142
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9968 6254 9996 8486
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 8294 10456 8434
rect 10520 8362 10548 9522
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9784 5370 9812 5578
rect 9954 5536 10010 5545
rect 9954 5471 10010 5480
rect 9862 5400 9918 5409
rect 9772 5364 9824 5370
rect 9862 5335 9918 5344
rect 9772 5306 9824 5312
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4078 9720 4966
rect 9784 4622 9812 5306
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9404 3936 9456 3942
rect 9402 3904 9404 3913
rect 9456 3904 9458 3913
rect 9402 3839 9458 3848
rect 9876 3738 9904 5335
rect 9968 5302 9996 5471
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 10060 4826 10088 7346
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10046 4720 10102 4729
rect 10046 4655 10102 4664
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9588 3528 9640 3534
rect 9640 3476 9720 3482
rect 9588 3470 9720 3476
rect 9600 3454 9720 3470
rect 9692 2825 9720 3454
rect 9678 2816 9734 2825
rect 9678 2751 9734 2760
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9968 2378 9996 2586
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9036 1896 9088 1902
rect 9036 1838 9088 1844
rect 8576 1828 8628 1834
rect 8576 1770 8628 1776
rect 9692 870 9812 898
rect 9692 800 9720 870
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 9784 762 9812 870
rect 10060 762 10088 4655
rect 10152 2650 10180 5646
rect 10244 3505 10272 8230
rect 10414 7848 10470 7857
rect 10414 7783 10470 7792
rect 10428 7410 10456 7783
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10336 4690 10364 6666
rect 10612 5846 10640 10678
rect 10704 7410 10732 11766
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 8945 10824 10406
rect 10874 9344 10930 9353
rect 10874 9279 10930 9288
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 10796 8498 10824 8871
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10416 5840 10468 5846
rect 10600 5840 10652 5846
rect 10416 5782 10468 5788
rect 10506 5808 10562 5817
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10230 3496 10286 3505
rect 10230 3431 10286 3440
rect 10244 3058 10272 3431
rect 10428 3194 10456 5782
rect 10600 5782 10652 5788
rect 10506 5743 10562 5752
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10520 2378 10548 5743
rect 10600 5704 10652 5710
rect 10796 5692 10824 8434
rect 10888 8430 10916 9279
rect 10980 9042 11008 15807
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 14006 11100 15370
rect 11256 15178 11284 18022
rect 11348 17202 11376 18958
rect 11426 18864 11482 18873
rect 11716 18850 11744 24618
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 11900 24410 11928 24550
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11794 22264 11850 22273
rect 11794 22199 11850 22208
rect 11808 22098 11836 22199
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11900 21894 11928 22034
rect 11888 21888 11940 21894
rect 11794 21856 11850 21865
rect 11888 21830 11940 21836
rect 11794 21791 11850 21800
rect 11426 18799 11482 18808
rect 11532 18822 11744 18850
rect 11440 18601 11468 18799
rect 11426 18592 11482 18601
rect 11426 18527 11482 18536
rect 11532 18358 11560 18822
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11716 18426 11744 18634
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11532 17746 11560 18158
rect 11520 17740 11572 17746
rect 11808 17728 11836 21791
rect 11888 21480 11940 21486
rect 11888 21422 11940 21428
rect 11900 18442 11928 21422
rect 11992 19768 12020 26726
rect 12268 26382 12296 27270
rect 12360 26994 12388 27474
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12452 25242 12480 29990
rect 13556 27470 13584 36722
rect 15396 34746 15424 36722
rect 15384 34740 15436 34746
rect 15384 34682 15436 34688
rect 13912 34604 13964 34610
rect 13912 34546 13964 34552
rect 13924 31754 13952 34546
rect 14188 31884 14240 31890
rect 14188 31826 14240 31832
rect 13832 31726 13952 31754
rect 13544 27464 13596 27470
rect 13544 27406 13596 27412
rect 13636 27464 13688 27470
rect 13636 27406 13688 27412
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12544 25362 12572 26726
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12072 25220 12124 25226
rect 12452 25214 12572 25242
rect 12072 25162 12124 25168
rect 12084 24954 12112 25162
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 12084 19922 12112 24890
rect 12544 24274 12572 25214
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12636 24138 12664 27270
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 12912 25498 12940 25842
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12716 24336 12768 24342
rect 12716 24278 12768 24284
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12452 23866 12480 24006
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12348 22500 12400 22506
rect 12348 22442 12400 22448
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12268 21622 12296 21830
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 12176 19786 12204 21286
rect 12360 21162 12388 22442
rect 12452 22030 12480 22918
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12268 21134 12388 21162
rect 12164 19780 12216 19786
rect 11992 19740 12112 19768
rect 12084 18873 12112 19740
rect 12164 19722 12216 19728
rect 12070 18864 12126 18873
rect 12070 18799 12126 18808
rect 12164 18760 12216 18766
rect 12162 18728 12164 18737
rect 12216 18728 12218 18737
rect 12162 18663 12218 18672
rect 11980 18624 12032 18630
rect 11978 18592 11980 18601
rect 12032 18592 12034 18601
rect 11978 18527 12034 18536
rect 11900 18414 12020 18442
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11900 17785 11928 18294
rect 11520 17682 11572 17688
rect 11716 17700 11836 17728
rect 11886 17776 11942 17785
rect 11886 17711 11942 17720
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11532 16998 11560 17682
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11348 15745 11376 16118
rect 11334 15736 11390 15745
rect 11334 15671 11390 15680
rect 11256 15150 11376 15178
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11150 14648 11206 14657
rect 11150 14583 11206 14592
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 11164 12764 11192 14583
rect 11256 13394 11284 14758
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11256 12918 11284 13126
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11072 12736 11192 12764
rect 11244 12776 11296 12782
rect 11072 10606 11100 12736
rect 11244 12718 11296 12724
rect 11152 12640 11204 12646
rect 11150 12608 11152 12617
rect 11204 12608 11206 12617
rect 11150 12543 11206 12552
rect 11256 12306 11284 12718
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11150 11928 11206 11937
rect 11150 11863 11206 11872
rect 11164 11694 11192 11863
rect 11256 11694 11284 12106
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11242 11112 11298 11121
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 11072 8820 11100 10066
rect 11164 9994 11192 11086
rect 11348 11082 11376 15150
rect 11440 13297 11468 16934
rect 11532 16658 11560 16934
rect 11624 16697 11652 17002
rect 11610 16688 11666 16697
rect 11520 16652 11572 16658
rect 11610 16623 11666 16632
rect 11520 16594 11572 16600
rect 11532 16046 11560 16594
rect 11716 16153 11744 17700
rect 11900 17610 11928 17711
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11992 17270 12020 18414
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12084 18057 12112 18294
rect 12070 18048 12126 18057
rect 12268 18034 12296 21134
rect 12544 20602 12572 23054
rect 12636 22710 12664 23462
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12728 22574 12756 24278
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 21486 12756 22510
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12636 20482 12664 21014
rect 12544 20454 12664 20482
rect 12438 19272 12494 19281
rect 12438 19207 12494 19216
rect 12452 18766 12480 19207
rect 12544 19174 12572 20454
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12636 19378 12664 20334
rect 12716 19712 12768 19718
rect 12714 19680 12716 19689
rect 12768 19680 12770 19689
rect 12714 19615 12770 19624
rect 12624 19372 12676 19378
rect 12676 19332 12756 19360
rect 12624 19314 12676 19320
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12360 18465 12388 18634
rect 12346 18456 12402 18465
rect 12346 18391 12402 18400
rect 12070 17983 12126 17992
rect 12176 18006 12296 18034
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 12084 17270 12112 17818
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 11992 16980 12020 17206
rect 11992 16952 12112 16980
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11702 16144 11758 16153
rect 11702 16079 11758 16088
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11532 14958 11560 15982
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11532 14482 11560 14894
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11624 14362 11652 15506
rect 11532 14334 11652 14362
rect 11426 13288 11482 13297
rect 11532 13258 11560 14334
rect 11716 14328 11744 16079
rect 11808 15706 11836 16730
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11796 14340 11848 14346
rect 11716 14300 11796 14328
rect 11796 14282 11848 14288
rect 11702 14240 11758 14249
rect 11702 14175 11758 14184
rect 11716 13938 11744 14175
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11716 13394 11744 13874
rect 11704 13388 11756 13394
rect 11900 13376 11928 16594
rect 12084 16538 12112 16952
rect 12176 16658 12204 18006
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12268 17746 12296 17818
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12360 16833 12388 17682
rect 12346 16824 12402 16833
rect 12346 16759 12402 16768
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12084 16510 12204 16538
rect 12070 16144 12126 16153
rect 12070 16079 12126 16088
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 14346 12020 15846
rect 12084 14958 12112 16079
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12084 14657 12112 14894
rect 12070 14648 12126 14657
rect 12070 14583 12126 14592
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11992 13530 12020 13806
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11900 13348 12020 13376
rect 11704 13330 11756 13336
rect 11426 13223 11482 13232
rect 11520 13252 11572 13258
rect 11440 12170 11468 13223
rect 11520 13194 11572 13200
rect 11532 12753 11560 13194
rect 11716 12850 11744 13330
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11518 12744 11574 12753
rect 11518 12679 11574 12688
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11716 11898 11744 12786
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11808 12073 11836 12106
rect 11794 12064 11850 12073
rect 11794 11999 11850 12008
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11242 11047 11298 11056
rect 11336 11076 11388 11082
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11164 9586 11192 9930
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10980 8792 11100 8820
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10888 6254 10916 8366
rect 10980 8129 11008 8792
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10966 8120 11022 8129
rect 11164 8072 11192 8434
rect 11256 8430 11284 11047
rect 11336 11018 11388 11024
rect 11334 10840 11390 10849
rect 11440 10826 11468 11698
rect 11390 10798 11468 10826
rect 11334 10775 11390 10784
rect 11348 10674 11376 10775
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 10966 8055 11022 8064
rect 10980 8022 11008 8055
rect 11072 8044 11192 8072
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11072 7886 11100 8044
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 7449 11008 7754
rect 11164 7721 11192 7890
rect 11150 7712 11206 7721
rect 11150 7647 11206 7656
rect 11150 7576 11206 7585
rect 11150 7511 11206 7520
rect 10966 7440 11022 7449
rect 10966 7375 11022 7384
rect 11058 7304 11114 7313
rect 11058 7239 11114 7248
rect 11072 6662 11100 7239
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10888 5846 10916 6054
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10652 5664 10824 5692
rect 10888 5681 10916 5782
rect 10874 5672 10930 5681
rect 10600 5646 10652 5652
rect 10612 2825 10640 5646
rect 10874 5607 10930 5616
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10704 3058 10732 4762
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10598 2816 10654 2825
rect 10598 2751 10654 2760
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 10796 1970 10824 5170
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10888 2106 10916 4150
rect 10980 4078 11008 4558
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 11072 2990 11100 6054
rect 11164 5098 11192 7511
rect 11256 7342 11284 8230
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11348 6662 11376 10134
rect 11532 9489 11560 11834
rect 11716 11762 11744 11834
rect 11992 11830 12020 13348
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12084 12345 12112 13194
rect 12176 13002 12204 16510
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12268 15502 12296 16118
rect 12360 15609 12388 16759
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12346 15600 12402 15609
rect 12346 15535 12402 15544
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12452 15366 12480 15642
rect 12544 15586 12572 19110
rect 12728 16726 12756 19332
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12544 15558 12756 15586
rect 12820 15570 12848 25298
rect 12912 25158 12940 25434
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12912 23338 12940 25094
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13188 24410 13216 24618
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23662 13032 24074
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 13096 23526 13124 24346
rect 13268 24336 13320 24342
rect 13268 24278 13320 24284
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 12912 23310 13124 23338
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12912 22030 12940 22374
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12912 21078 12940 21966
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 12912 19310 12940 20266
rect 13004 19310 13032 21354
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 13004 18329 13032 18362
rect 12990 18320 13046 18329
rect 12990 18255 13046 18264
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 12912 16250 12940 16662
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12544 15201 12572 15438
rect 12254 15192 12310 15201
rect 12254 15127 12310 15136
rect 12530 15192 12586 15201
rect 12530 15127 12586 15136
rect 12268 14770 12296 15127
rect 12268 14742 12388 14770
rect 12360 13190 12388 14742
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12176 12974 12388 13002
rect 12070 12336 12126 12345
rect 12070 12271 12126 12280
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11992 11218 12020 11766
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11900 10810 11928 11018
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 12072 10600 12124 10606
rect 12176 10554 12204 10746
rect 12268 10742 12296 12106
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12360 10606 12388 12974
rect 12452 12434 12480 13942
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12782 12664 13330
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12728 12442 12756 15558
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12912 15162 12940 15370
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13004 12458 13032 16594
rect 13096 13326 13124 23310
rect 13188 22710 13216 24210
rect 13280 23186 13308 24278
rect 13372 23497 13400 24550
rect 13358 23488 13414 23497
rect 13358 23423 13414 23432
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 13188 21010 13216 22646
rect 13358 22264 13414 22273
rect 13358 22199 13414 22208
rect 13268 22024 13320 22030
rect 13266 21992 13268 22001
rect 13320 21992 13322 22001
rect 13266 21927 13322 21936
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13280 21078 13308 21422
rect 13268 21072 13320 21078
rect 13268 21014 13320 21020
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13372 20924 13400 22199
rect 13280 20896 13400 20924
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13188 19990 13216 20470
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13176 19780 13228 19786
rect 13176 19722 13228 19728
rect 13188 19242 13216 19722
rect 13176 19236 13228 19242
rect 13176 19178 13228 19184
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13188 16794 13216 17546
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13280 16674 13308 20896
rect 13358 20360 13414 20369
rect 13464 20330 13492 27270
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13556 24274 13584 24550
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13648 22094 13676 27406
rect 13832 26858 13860 31726
rect 14200 27878 14228 31826
rect 15580 28558 15608 37062
rect 16776 36922 16804 39200
rect 17420 37126 17448 39200
rect 17500 37256 17552 37262
rect 17500 37198 17552 37204
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 16764 36916 16816 36922
rect 16764 36858 16816 36864
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17132 30592 17184 30598
rect 17132 30534 17184 30540
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15200 28144 15252 28150
rect 15200 28086 15252 28092
rect 14188 27872 14240 27878
rect 14188 27814 14240 27820
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14384 27062 14412 27270
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14476 26994 14504 27338
rect 15212 27130 15240 28086
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 13820 26852 13872 26858
rect 13820 26794 13872 26800
rect 13912 26852 13964 26858
rect 13912 26794 13964 26800
rect 13924 26450 13952 26794
rect 13912 26444 13964 26450
rect 13912 26386 13964 26392
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13740 23798 13768 25230
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13832 24274 13860 24754
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13728 23792 13780 23798
rect 13728 23734 13780 23740
rect 13740 23662 13768 23734
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13924 23594 13952 26386
rect 14016 26042 14044 26862
rect 14004 26036 14056 26042
rect 14004 25978 14056 25984
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 14108 24886 14136 25638
rect 14924 25356 14976 25362
rect 14924 25298 14976 25304
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 14372 24744 14424 24750
rect 14424 24692 14688 24698
rect 14372 24686 14688 24692
rect 14384 24682 14688 24686
rect 14384 24676 14700 24682
rect 14384 24670 14648 24676
rect 14648 24618 14700 24624
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 14384 23254 14412 24006
rect 14830 23760 14886 23769
rect 14830 23695 14832 23704
rect 14884 23695 14886 23704
rect 14832 23666 14884 23672
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13832 22710 13860 23122
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14108 22710 14136 22918
rect 14292 22778 14320 22918
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 13648 22066 13768 22094
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13648 21010 13676 21354
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13648 20602 13676 20810
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13358 20295 13414 20304
rect 13452 20324 13504 20330
rect 13188 16646 13308 16674
rect 13372 16658 13400 20295
rect 13452 20266 13504 20272
rect 13556 19922 13584 20470
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13740 19334 13768 22066
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14186 21584 14242 21593
rect 14186 21519 14188 21528
rect 14240 21519 14242 21528
rect 14188 21490 14240 21496
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13648 19306 13768 19334
rect 13450 18592 13506 18601
rect 13450 18527 13506 18536
rect 13464 18358 13492 18527
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13450 18184 13506 18193
rect 13450 18119 13506 18128
rect 13464 18086 13492 18119
rect 13556 18086 13584 19246
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13648 17490 13676 19306
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13556 17462 13676 17490
rect 13360 16652 13412 16658
rect 13188 15570 13216 16646
rect 13360 16594 13412 16600
rect 13358 16280 13414 16289
rect 13268 16244 13320 16250
rect 13358 16215 13414 16224
rect 13268 16186 13320 16192
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13174 12744 13230 12753
rect 13174 12679 13230 12688
rect 12716 12436 12768 12442
rect 12452 12406 12572 12434
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12452 11014 12480 11766
rect 12544 11558 12572 12406
rect 13004 12430 13124 12458
rect 12716 12378 12768 12384
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12912 11286 12940 12106
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12124 10548 12204 10554
rect 12072 10542 12204 10548
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 11610 10024 11666 10033
rect 11610 9959 11666 9968
rect 11518 9480 11574 9489
rect 11518 9415 11574 9424
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11532 8945 11560 9114
rect 11624 9042 11652 9959
rect 11716 9450 11744 10542
rect 12084 10526 12204 10542
rect 11888 10192 11940 10198
rect 11886 10160 11888 10169
rect 11940 10160 11942 10169
rect 11886 10095 11942 10104
rect 12162 10024 12218 10033
rect 12162 9959 12164 9968
rect 12216 9959 12218 9968
rect 12808 9988 12860 9994
rect 12164 9930 12216 9936
rect 12808 9930 12860 9936
rect 11796 9512 11848 9518
rect 12164 9512 12216 9518
rect 11848 9472 11928 9500
rect 11796 9454 11848 9460
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11518 8936 11574 8945
rect 11518 8871 11574 8880
rect 11716 8498 11744 9386
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11808 9217 11836 9318
rect 11794 9208 11850 9217
rect 11794 9143 11850 9152
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11900 8106 11928 9472
rect 12164 9454 12216 9460
rect 12176 8265 12204 9454
rect 12530 9208 12586 9217
rect 12530 9143 12586 9152
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8566 12388 8910
rect 12544 8838 12572 9143
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12162 8256 12218 8265
rect 12162 8191 12218 8200
rect 11900 8078 12204 8106
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7426 11744 7890
rect 12070 7712 12126 7721
rect 12070 7647 12126 7656
rect 12084 7478 12112 7647
rect 11532 7398 11744 7426
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11256 5778 11284 6190
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11256 5234 11284 5714
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11164 4321 11192 5034
rect 11440 4554 11468 6326
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11150 4312 11206 4321
rect 11150 4247 11206 4256
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11256 2922 11284 3334
rect 11440 2990 11468 4490
rect 11532 3913 11560 7398
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11624 6254 11652 7278
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11900 6458 11928 6598
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11624 5778 11652 6190
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11900 5574 11928 5850
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 12070 5264 12126 5273
rect 12070 5199 12126 5208
rect 11704 5160 11756 5166
rect 11978 5128 12034 5137
rect 11756 5108 11836 5114
rect 11704 5102 11836 5108
rect 11716 5086 11836 5102
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11612 3936 11664 3942
rect 11518 3904 11574 3913
rect 11612 3878 11664 3884
rect 11518 3839 11574 3848
rect 11624 3670 11652 3878
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11716 2514 11744 4014
rect 11808 3602 11836 5086
rect 11978 5063 12034 5072
rect 11992 4690 12020 5063
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 12084 4457 12112 5199
rect 12176 5114 12204 8078
rect 12360 7534 12572 7562
rect 12360 6338 12388 7534
rect 12544 7460 12572 7534
rect 12624 7472 12676 7478
rect 12544 7432 12624 7460
rect 12624 7414 12676 7420
rect 12728 7324 12756 8366
rect 12268 6310 12388 6338
rect 12544 7296 12756 7324
rect 12268 5545 12296 6310
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12254 5536 12310 5545
rect 12254 5471 12310 5480
rect 12360 5273 12388 6190
rect 12346 5264 12402 5273
rect 12346 5199 12402 5208
rect 12176 5086 12296 5114
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12176 4593 12204 4966
rect 12162 4584 12218 4593
rect 12162 4519 12218 4528
rect 12070 4448 12126 4457
rect 12070 4383 12126 4392
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 12162 3904 12218 3913
rect 11992 3738 12020 3878
rect 12162 3839 12218 3848
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11808 3058 11836 3538
rect 11980 3528 12032 3534
rect 11978 3496 11980 3505
rect 12032 3496 12034 3505
rect 12176 3466 12204 3839
rect 12268 3738 12296 5086
rect 12544 4826 12572 7296
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12622 6080 12678 6089
rect 12622 6015 12678 6024
rect 12636 5681 12664 6015
rect 12622 5672 12678 5681
rect 12622 5607 12678 5616
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12346 4448 12402 4457
rect 12346 4383 12402 4392
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12360 3602 12388 4383
rect 12452 3942 12480 4694
rect 12530 4584 12586 4593
rect 12530 4519 12586 4528
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 11978 3431 12034 3440
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 12544 2774 12572 4519
rect 12728 2854 12756 6666
rect 12820 3194 12848 9930
rect 12912 7206 12940 11086
rect 13096 10985 13124 12430
rect 13082 10976 13138 10985
rect 13082 10911 13138 10920
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6730 12940 7142
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12898 6488 12954 6497
rect 12898 6423 12954 6432
rect 12912 4826 12940 6423
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12544 2746 12664 2774
rect 12636 2650 12664 2746
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 9784 734 10088 762
rect 10888 870 11008 898
rect 10888 202 10916 870
rect 10980 800 11008 870
rect 11624 870 11744 898
rect 11624 800 11652 870
rect 10876 196 10928 202
rect 10966 200 11022 800
rect 11610 200 11666 800
rect 10876 138 10928 144
rect 11716 134 11744 870
rect 12912 800 12940 4218
rect 13004 2774 13032 8502
rect 13096 6474 13124 9862
rect 13188 9450 13216 12679
rect 13280 10742 13308 16186
rect 13372 16046 13400 16215
rect 13360 16040 13412 16046
rect 13412 16000 13492 16028
rect 13360 15982 13412 15988
rect 13360 15904 13412 15910
rect 13358 15872 13360 15881
rect 13412 15872 13414 15881
rect 13358 15807 13414 15816
rect 13358 15600 13414 15609
rect 13358 15535 13414 15544
rect 13372 15162 13400 15535
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13464 14074 13492 16000
rect 13556 15638 13584 17462
rect 13634 17368 13690 17377
rect 13634 17303 13690 17312
rect 13648 17202 13676 17303
rect 13740 17241 13768 19110
rect 13832 18465 13860 19926
rect 14002 19408 14058 19417
rect 14002 19343 14058 19352
rect 13818 18456 13874 18465
rect 13818 18391 13874 18400
rect 13820 17536 13872 17542
rect 13818 17504 13820 17513
rect 13872 17504 13874 17513
rect 13874 17462 13952 17490
rect 13818 17439 13874 17448
rect 13726 17232 13782 17241
rect 13636 17196 13688 17202
rect 13726 17167 13782 17176
rect 13636 17138 13688 17144
rect 13818 16688 13874 16697
rect 13818 16623 13874 16632
rect 13832 16046 13860 16623
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12617 13492 13262
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13450 12608 13506 12617
rect 13450 12543 13506 12552
rect 13556 12442 13584 13194
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8809 13308 8910
rect 13266 8800 13322 8809
rect 13266 8735 13322 8744
rect 13268 8628 13320 8634
rect 13372 8616 13400 12174
rect 13648 11937 13676 13398
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12918 13768 13126
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13634 11928 13690 11937
rect 13634 11863 13690 11872
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11218 13492 11494
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 10198 13492 11154
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13648 9674 13676 11863
rect 13740 11286 13768 12378
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13740 10470 13768 11018
rect 13832 10849 13860 14758
rect 13924 14550 13952 17462
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 14016 14090 14044 19343
rect 14108 19258 14136 21014
rect 14292 20856 14320 21830
rect 14384 21350 14412 22510
rect 14752 22094 14780 23258
rect 14844 23254 14872 23666
rect 14832 23248 14884 23254
rect 14832 23190 14884 23196
rect 14936 23202 14964 25298
rect 15108 24812 15160 24818
rect 15108 24754 15160 24760
rect 15120 24206 15148 24754
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15016 24064 15068 24070
rect 15016 24006 15068 24012
rect 15028 23866 15056 24006
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 15120 23322 15148 23802
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 14936 23174 15148 23202
rect 15212 23186 15240 24550
rect 15660 23588 15712 23594
rect 15660 23530 15712 23536
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 14752 22066 14872 22094
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14476 21622 14504 21830
rect 14464 21616 14516 21622
rect 14464 21558 14516 21564
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14384 21078 14412 21286
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14568 20874 14596 21898
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14556 20868 14608 20874
rect 14292 20828 14504 20856
rect 14370 20360 14426 20369
rect 14370 20295 14426 20304
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14200 19446 14228 19654
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14108 19230 14228 19258
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14108 16590 14136 18702
rect 14200 18698 14228 19230
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14200 18601 14228 18634
rect 14280 18624 14332 18630
rect 14186 18592 14242 18601
rect 14280 18566 14332 18572
rect 14186 18527 14242 18536
rect 14292 18358 14320 18566
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14188 17604 14240 17610
rect 14188 17546 14240 17552
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14108 16425 14136 16526
rect 14094 16416 14150 16425
rect 14094 16351 14150 16360
rect 13924 14062 14044 14090
rect 13924 13734 13952 14062
rect 14096 14000 14148 14006
rect 14200 13988 14228 17546
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14292 15881 14320 16050
rect 14278 15872 14334 15881
rect 14278 15807 14334 15816
rect 14280 14000 14332 14006
rect 14200 13960 14280 13988
rect 14096 13942 14148 13948
rect 14280 13942 14332 13948
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14016 12238 14044 12718
rect 14108 12714 14136 13942
rect 14278 13696 14334 13705
rect 14278 13631 14334 13640
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13818 10840 13874 10849
rect 13818 10775 13874 10784
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13556 9646 13676 9674
rect 13556 9602 13584 9646
rect 13320 8588 13400 8616
rect 13268 8570 13320 8576
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13188 7426 13216 7482
rect 13188 7398 13308 7426
rect 13096 6446 13216 6474
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13096 5914 13124 6258
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13188 3738 13216 6446
rect 13280 5953 13308 7398
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6118 13400 6598
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13266 5944 13322 5953
rect 13266 5879 13322 5888
rect 13280 5846 13308 5879
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13266 5672 13322 5681
rect 13266 5607 13322 5616
rect 13280 4078 13308 5607
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13372 3398 13400 4966
rect 13464 4826 13492 9590
rect 13556 9574 13676 9602
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13556 8090 13584 8502
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13648 7954 13676 9574
rect 13740 8974 13768 9930
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 13556 5817 13584 6151
rect 13542 5808 13598 5817
rect 13542 5743 13598 5752
rect 13556 5710 13584 5743
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13542 4448 13598 4457
rect 13542 4383 13598 4392
rect 13450 4040 13506 4049
rect 13450 3975 13506 3984
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13464 3194 13492 3975
rect 13556 3670 13584 4383
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13740 2990 13768 8298
rect 13832 7478 13860 10775
rect 13924 8634 13952 12038
rect 14016 11898 14044 12174
rect 14108 12073 14136 12242
rect 14094 12064 14150 12073
rect 14094 11999 14150 12008
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14016 10606 14044 11086
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 9518 14044 10542
rect 14200 9654 14228 12854
rect 14292 12753 14320 13631
rect 14384 13394 14412 20295
rect 14476 19786 14504 20828
rect 14556 20810 14608 20816
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14462 19680 14518 19689
rect 14462 19615 14518 19624
rect 14476 18222 14504 19615
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14568 18698 14596 18770
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14554 18320 14610 18329
rect 14554 18255 14610 18264
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14476 17338 14504 17546
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14568 15978 14596 18255
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14476 13530 14504 14350
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14278 12744 14334 12753
rect 14278 12679 14334 12688
rect 14292 12434 14320 12679
rect 14292 12406 14412 12434
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 10169 14320 10542
rect 14278 10160 14334 10169
rect 14278 10095 14334 10104
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14292 9042 14320 9454
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14004 8968 14056 8974
rect 14056 8928 14136 8956
rect 14004 8910 14056 8916
rect 14108 8673 14136 8928
rect 14186 8800 14242 8809
rect 14186 8735 14242 8744
rect 14094 8664 14150 8673
rect 13912 8628 13964 8634
rect 14094 8599 14150 8608
rect 13912 8570 13964 8576
rect 14108 8430 14136 8599
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14200 8090 14228 8735
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14002 7848 14058 7857
rect 14002 7783 14058 7792
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 14016 6866 14044 7783
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 4282 13860 6666
rect 13910 5536 13966 5545
rect 13910 5471 13966 5480
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13924 4049 13952 5471
rect 14108 5001 14136 7482
rect 14200 7410 14228 8026
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 6866 14228 7346
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6633 14320 6734
rect 14278 6624 14334 6633
rect 14278 6559 14334 6568
rect 14094 4992 14150 5001
rect 14094 4927 14150 4936
rect 14002 4856 14058 4865
rect 14002 4791 14058 4800
rect 14016 4214 14044 4791
rect 14108 4622 14136 4927
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14200 4146 14228 4626
rect 14278 4584 14334 4593
rect 14278 4519 14280 4528
rect 14332 4519 14334 4528
rect 14280 4490 14332 4496
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14096 4072 14148 4078
rect 13910 4040 13966 4049
rect 13820 4004 13872 4010
rect 14096 4014 14148 4020
rect 13910 3975 13966 3984
rect 13820 3946 13872 3952
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13004 2746 13124 2774
rect 13096 2310 13124 2746
rect 13556 2514 13584 2926
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13740 1766 13768 2586
rect 13728 1760 13780 1766
rect 13728 1702 13780 1708
rect 13832 1630 13860 3946
rect 14108 1737 14136 4014
rect 14186 3768 14242 3777
rect 14186 3703 14242 3712
rect 14094 1728 14150 1737
rect 14094 1663 14150 1672
rect 13820 1624 13872 1630
rect 13820 1566 13872 1572
rect 14200 800 14228 3703
rect 14280 3664 14332 3670
rect 14384 3641 14412 12406
rect 14476 11200 14504 13466
rect 14568 12628 14596 15914
rect 14660 13870 14688 20946
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14752 17134 14780 20810
rect 14844 17542 14872 22066
rect 14922 21992 14978 22001
rect 14922 21927 14978 21936
rect 14936 21554 14964 21927
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14936 19514 14964 21490
rect 15028 21010 15056 22170
rect 15120 22098 15148 23174
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15488 22778 15516 23462
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 15212 21962 15240 22374
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15200 20936 15252 20942
rect 15028 20884 15200 20890
rect 15028 20878 15252 20884
rect 15028 20862 15240 20878
rect 15028 20505 15056 20862
rect 15200 20800 15252 20806
rect 15304 20777 15332 22102
rect 15396 20806 15424 22170
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15384 20800 15436 20806
rect 15200 20742 15252 20748
rect 15290 20768 15346 20777
rect 15014 20496 15070 20505
rect 15014 20431 15070 20440
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15120 19514 15148 20402
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14844 16182 14872 16458
rect 14832 16176 14884 16182
rect 14832 16118 14884 16124
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15706 14780 16050
rect 14740 15700 14792 15706
rect 14936 15688 14964 18362
rect 15028 18290 15056 18362
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15014 18184 15070 18193
rect 15014 18119 15016 18128
rect 15068 18119 15070 18128
rect 15016 18090 15068 18096
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 15028 16522 15056 17682
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14740 15642 14792 15648
rect 14844 15660 14964 15688
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14752 12986 14780 15642
rect 14844 15366 14872 15660
rect 15028 15620 15056 16458
rect 14936 15592 15056 15620
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14936 13025 14964 15592
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 15094 15056 15370
rect 15016 15088 15068 15094
rect 15014 15056 15016 15065
rect 15068 15056 15070 15065
rect 15014 14991 15070 15000
rect 15120 14550 15148 19314
rect 15212 17270 15240 20742
rect 15384 20742 15436 20748
rect 15290 20703 15346 20712
rect 15488 20534 15516 21286
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15396 19786 15424 19994
rect 15474 19816 15530 19825
rect 15384 19780 15436 19786
rect 15436 19760 15474 19768
rect 15436 19751 15530 19760
rect 15436 19740 15516 19751
rect 15384 19722 15436 19728
rect 15382 19544 15438 19553
rect 15382 19479 15438 19488
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15304 17785 15332 19178
rect 15290 17776 15346 17785
rect 15290 17711 15346 17720
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15304 16289 15332 17614
rect 15396 17610 15424 19479
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15396 17513 15424 17546
rect 15382 17504 15438 17513
rect 15382 17439 15438 17448
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15290 16280 15346 16289
rect 15290 16215 15346 16224
rect 15396 15978 15424 16934
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15212 14482 15240 15438
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15304 14822 15332 15370
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15396 14634 15424 15914
rect 15488 15314 15516 19740
rect 15580 18970 15608 22986
rect 15672 22982 15700 23530
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15672 20398 15700 22918
rect 15764 22234 15792 28358
rect 16396 26308 16448 26314
rect 16396 26250 16448 26256
rect 15936 25764 15988 25770
rect 15936 25706 15988 25712
rect 15948 23730 15976 25706
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 16224 24410 16252 24618
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15934 22264 15990 22273
rect 15752 22228 15804 22234
rect 15934 22199 15990 22208
rect 15752 22170 15804 22176
rect 15948 22098 15976 22199
rect 16040 22137 16068 22578
rect 16026 22128 16082 22137
rect 15936 22092 15988 22098
rect 16026 22063 16082 22072
rect 15936 22034 15988 22040
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16132 21146 16160 21422
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 15844 21072 15896 21078
rect 16028 21072 16080 21078
rect 15896 21020 16028 21026
rect 15844 21014 16080 21020
rect 15856 20998 16068 21014
rect 16224 20942 16252 21082
rect 16212 20936 16264 20942
rect 15764 20874 15976 20890
rect 16212 20878 16264 20884
rect 15764 20868 15988 20874
rect 15764 20862 15936 20868
rect 15764 20806 15792 20862
rect 15936 20810 15988 20816
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15842 20496 15898 20505
rect 15842 20431 15898 20440
rect 15660 20392 15712 20398
rect 15658 20360 15660 20369
rect 15712 20360 15714 20369
rect 15658 20295 15714 20304
rect 15658 19952 15714 19961
rect 15658 19887 15714 19896
rect 15672 19378 15700 19887
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 16114 15608 16526
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15566 15736 15622 15745
rect 15566 15671 15622 15680
rect 15580 15638 15608 15671
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15488 15286 15608 15314
rect 15474 15192 15530 15201
rect 15474 15127 15530 15136
rect 15304 14606 15424 14634
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14922 13016 14978 13025
rect 14740 12980 14792 12986
rect 14922 12951 14978 12960
rect 14740 12922 14792 12928
rect 15028 12646 15056 14010
rect 15212 14006 15240 14418
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15120 13190 15148 13670
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15016 12640 15068 12646
rect 14568 12600 14964 12628
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14568 11830 14596 12242
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14556 11212 14608 11218
rect 14476 11172 14556 11200
rect 14556 11154 14608 11160
rect 14660 11098 14688 11834
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14568 11082 14688 11098
rect 14556 11076 14688 11082
rect 14608 11070 14688 11076
rect 14556 11018 14608 11024
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 8498 14504 9318
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14568 8129 14596 8842
rect 14752 8786 14780 11766
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14844 10606 14872 10950
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14660 8758 14780 8786
rect 14554 8120 14610 8129
rect 14554 8055 14610 8064
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 5930 14596 7686
rect 14660 6905 14688 8758
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14646 6896 14702 6905
rect 14752 6866 14780 8502
rect 14646 6831 14702 6840
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14568 5902 14780 5930
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14280 3606 14332 3612
rect 14370 3632 14426 3641
rect 14292 3466 14320 3606
rect 14370 3567 14426 3576
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14476 2961 14504 5578
rect 14660 5302 14688 5714
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14660 4690 14688 5238
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14556 4548 14608 4554
rect 14556 4490 14608 4496
rect 14568 4078 14596 4490
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14568 3466 14596 3674
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14752 3398 14780 5902
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14462 2952 14518 2961
rect 14462 2887 14518 2896
rect 14844 2650 14872 10406
rect 14936 10130 14964 12600
rect 15120 12617 15148 12922
rect 15016 12582 15068 12588
rect 15106 12608 15162 12617
rect 15106 12543 15162 12552
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 14936 7342 14964 8978
rect 15028 8945 15056 12106
rect 15014 8936 15070 8945
rect 15014 8871 15070 8880
rect 15120 8566 15148 12543
rect 15198 12064 15254 12073
rect 15198 11999 15254 12008
rect 15212 9722 15240 11999
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15120 8430 15148 8502
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15212 8294 15240 8842
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14922 6488 14978 6497
rect 14922 6423 14978 6432
rect 14936 6390 14964 6423
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14936 4486 14964 4762
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15028 3913 15056 5578
rect 15014 3904 15070 3913
rect 15014 3839 15070 3848
rect 15120 3194 15148 6666
rect 15212 6662 15240 7890
rect 15304 7342 15332 14606
rect 15488 14482 15516 15127
rect 15580 14958 15608 15286
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15384 13388 15436 13394
rect 15488 13376 15516 13806
rect 15436 13348 15516 13376
rect 15384 13330 15436 13336
rect 15396 9518 15424 13330
rect 15474 11384 15530 11393
rect 15474 11319 15530 11328
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15488 7585 15516 11319
rect 15580 10130 15608 14418
rect 15764 13433 15792 19790
rect 15856 19242 15884 20431
rect 16408 20058 16436 26250
rect 17144 25362 17172 30534
rect 17224 30116 17276 30122
rect 17224 30058 17276 30064
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16960 24750 16988 25094
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 17052 23526 17080 24550
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16592 21049 16620 22510
rect 16776 22166 16804 22918
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 16578 21040 16634 21049
rect 16578 20975 16634 20984
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16684 19718 16712 19858
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15856 16794 15884 17818
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15856 16114 15884 16458
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 15750 13424 15806 13433
rect 15750 13359 15806 13368
rect 15660 12776 15712 12782
rect 15658 12744 15660 12753
rect 15712 12744 15714 12753
rect 15658 12679 15714 12688
rect 15764 11558 15792 13359
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15856 10962 15884 15370
rect 15764 10934 15884 10962
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15580 8430 15608 10066
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15474 7576 15530 7585
rect 15474 7511 15530 7520
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15212 6254 15240 6598
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15304 5681 15332 6802
rect 15290 5672 15346 5681
rect 15290 5607 15346 5616
rect 15396 5409 15424 7414
rect 15382 5400 15438 5409
rect 15382 5335 15438 5344
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15212 3369 15240 3402
rect 15198 3360 15254 3369
rect 15198 3295 15254 3304
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14936 2825 14964 3062
rect 15304 2854 15332 4966
rect 15382 4176 15438 4185
rect 15382 4111 15438 4120
rect 15396 3194 15424 4111
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15672 2854 15700 10678
rect 15764 9382 15792 10934
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 9217 15792 9318
rect 15750 9208 15806 9217
rect 15750 9143 15806 9152
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15764 4185 15792 8366
rect 15856 5166 15884 10134
rect 15948 9926 15976 18022
rect 16040 12374 16068 18702
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16118 16824 16174 16833
rect 16118 16759 16120 16768
rect 16172 16759 16174 16768
rect 16120 16730 16172 16736
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 14929 16160 15438
rect 16118 14920 16174 14929
rect 16118 14855 16174 14864
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16132 13326 16160 13670
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 13025 16160 13262
rect 16118 13016 16174 13025
rect 16118 12951 16174 12960
rect 16028 12368 16080 12374
rect 16026 12336 16028 12345
rect 16080 12336 16082 12345
rect 16026 12271 16082 12280
rect 16224 12170 16252 18022
rect 16408 17066 16436 18702
rect 16592 17882 16620 19382
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16316 11286 16344 16050
rect 16408 12238 16436 17002
rect 16592 16969 16620 17478
rect 16578 16960 16634 16969
rect 16578 16895 16634 16904
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16592 15706 16620 15982
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16684 13394 16712 19654
rect 16776 18834 16804 22102
rect 17052 22098 17080 23462
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17144 21622 17172 22986
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16776 16658 16804 18770
rect 16868 18057 16896 21286
rect 17236 21010 17264 30058
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17328 23050 17356 26250
rect 17420 23186 17448 31962
rect 17512 31754 17540 37198
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 17776 32768 17828 32774
rect 17776 32710 17828 32716
rect 17512 31726 17724 31754
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17512 24954 17540 25298
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 17604 24154 17632 26318
rect 17512 24126 17632 24154
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17328 22953 17356 22986
rect 17314 22944 17370 22953
rect 17314 22879 17370 22888
rect 17512 21321 17540 24126
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17604 23798 17632 24006
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17696 23322 17724 31726
rect 17788 24410 17816 32710
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17776 24404 17828 24410
rect 17776 24346 17828 24352
rect 17880 24274 17908 25434
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17788 23798 17816 24210
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 17972 23662 18000 27882
rect 18064 26586 18092 36722
rect 18604 36372 18656 36378
rect 18604 36314 18656 36320
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18144 27872 18196 27878
rect 18144 27814 18196 27820
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 18156 24818 18184 27814
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18052 24336 18104 24342
rect 18052 24278 18104 24284
rect 18064 23866 18092 24278
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 18248 23594 18276 29990
rect 18616 26042 18644 36314
rect 18708 35834 18736 39200
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 18788 37188 18840 37194
rect 18788 37130 18840 37136
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 18800 25974 18828 37130
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19156 36848 19208 36854
rect 19156 36790 19208 36796
rect 19168 33522 19196 36790
rect 19156 33516 19208 33522
rect 19156 33458 19208 33464
rect 19168 28082 19196 33458
rect 19352 31822 19380 37062
rect 19444 35834 19472 37198
rect 19996 37126 20024 39200
rect 21284 37330 21312 39200
rect 21272 37324 21324 37330
rect 21272 37266 21324 37272
rect 20076 37256 20128 37262
rect 21928 37244 21956 39200
rect 21928 37216 22140 37244
rect 20076 37198 20128 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19064 26512 19116 26518
rect 19064 26454 19116 26460
rect 18788 25968 18840 25974
rect 18788 25910 18840 25916
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18800 25498 18828 25638
rect 18788 25492 18840 25498
rect 18788 25434 18840 25440
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18236 23588 18288 23594
rect 18236 23530 18288 23536
rect 17774 23488 17830 23497
rect 17774 23423 17830 23432
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17498 21312 17554 21321
rect 17498 21247 17554 21256
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 16960 20466 16988 20946
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16960 18222 16988 20402
rect 17130 20088 17186 20097
rect 17130 20023 17186 20032
rect 17144 19990 17172 20023
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17236 18970 17264 20470
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 17328 19922 17356 20198
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16854 18048 16910 18057
rect 16854 17983 16910 17992
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17236 17270 17264 17478
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16776 14618 16804 16458
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 15934 9480 15990 9489
rect 15934 9415 15990 9424
rect 15948 9382 15976 9415
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15948 5642 15976 8774
rect 16040 8022 16068 9590
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16132 6769 16160 9454
rect 16224 8974 16252 9998
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16316 8786 16344 11222
rect 16500 10538 16528 12038
rect 16592 11218 16620 12310
rect 16868 12306 16896 16934
rect 17052 16726 17080 17002
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17328 15502 17356 16118
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17040 15360 17092 15366
rect 17132 15360 17184 15366
rect 17040 15302 17092 15308
rect 17130 15328 17132 15337
rect 17184 15328 17186 15337
rect 17052 15094 17080 15302
rect 17130 15263 17186 15272
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 14006 17080 14214
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16684 11529 16712 12106
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16776 11898 16804 12038
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16960 11812 16988 13330
rect 17052 13297 17080 13330
rect 17038 13288 17094 13297
rect 17038 13223 17094 13232
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17038 12744 17094 12753
rect 17038 12679 17094 12688
rect 16868 11784 16988 11812
rect 16670 11520 16726 11529
rect 16670 11455 16726 11464
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16592 10266 16620 11154
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16408 9994 16436 10202
rect 16578 10160 16634 10169
rect 16578 10095 16634 10104
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16224 8758 16344 8786
rect 16118 6760 16174 6769
rect 16118 6695 16174 6704
rect 16132 6225 16160 6695
rect 16118 6216 16174 6225
rect 16118 6151 16174 6160
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 16028 5568 16080 5574
rect 16026 5536 16028 5545
rect 16120 5568 16172 5574
rect 16080 5536 16082 5545
rect 16120 5510 16172 5516
rect 16026 5471 16082 5480
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15948 4486 15976 5034
rect 15936 4480 15988 4486
rect 16040 4457 16068 5471
rect 15936 4422 15988 4428
rect 16026 4448 16082 4457
rect 15750 4176 15806 4185
rect 15750 4111 15806 4120
rect 15842 3632 15898 3641
rect 15842 3567 15898 3576
rect 15856 3466 15884 3567
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15948 3346 15976 4422
rect 16026 4383 16082 4392
rect 16132 3602 16160 5510
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15856 3318 15976 3346
rect 15292 2848 15344 2854
rect 14922 2816 14978 2825
rect 15292 2790 15344 2796
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 14922 2751 14978 2760
rect 15382 2680 15438 2689
rect 14832 2644 14884 2650
rect 15382 2615 15438 2624
rect 14832 2586 14884 2592
rect 15396 2446 15424 2615
rect 15856 2582 15884 3318
rect 16026 3224 16082 3233
rect 16026 3159 16028 3168
rect 16080 3159 16082 3168
rect 16028 3130 16080 3136
rect 16224 2972 16252 8758
rect 16408 8090 16436 9386
rect 16500 9110 16528 9522
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16592 8906 16620 10095
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16500 7886 16528 8230
rect 16578 8120 16634 8129
rect 16578 8055 16634 8064
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16592 7750 16620 8055
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16408 7262 16620 7290
rect 16408 7206 16436 7262
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 6866 16528 7142
rect 16592 7041 16620 7262
rect 16578 7032 16634 7041
rect 16578 6967 16634 6976
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16302 6760 16358 6769
rect 16302 6695 16358 6704
rect 16316 6322 16344 6695
rect 16304 6316 16356 6322
rect 16356 6276 16436 6304
rect 16304 6258 16356 6264
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16040 2944 16252 2972
rect 16040 2774 16068 2944
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15948 2746 16068 2774
rect 15844 2576 15896 2582
rect 15844 2518 15896 2524
rect 15948 2446 15976 2746
rect 16132 2650 16160 2790
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16316 2446 16344 3878
rect 16408 3369 16436 6276
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16500 5953 16528 6190
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16486 5944 16542 5953
rect 16486 5879 16542 5888
rect 16592 5817 16620 6054
rect 16578 5808 16634 5817
rect 16578 5743 16634 5752
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 4622 16620 5034
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16486 3632 16542 3641
rect 16486 3567 16542 3576
rect 16394 3360 16450 3369
rect 16394 3295 16450 3304
rect 16408 3194 16436 3295
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16500 3126 16528 3567
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16684 2904 16712 9998
rect 16776 8498 16804 10610
rect 16868 10198 16896 11784
rect 17052 11694 17080 12679
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 16960 10606 16988 11630
rect 17144 11626 17172 12922
rect 17236 12850 17264 13738
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17236 12170 17264 12650
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17236 11558 17264 12106
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17052 11286 17080 11494
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 17222 11248 17278 11257
rect 17222 11183 17278 11192
rect 17236 11082 17264 11183
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17038 10704 17094 10713
rect 17328 10674 17356 12582
rect 17038 10639 17094 10648
rect 17316 10668 17368 10674
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16762 6896 16818 6905
rect 16762 6831 16818 6840
rect 16776 5710 16804 6831
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 5234 16804 5510
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16868 5030 16896 9386
rect 16960 6254 16988 10542
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 17052 5114 17080 10639
rect 17316 10610 17368 10616
rect 17420 10130 17448 20946
rect 17512 19854 17540 21247
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17512 15978 17540 17546
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17604 15065 17632 22510
rect 17788 22094 17816 23423
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17696 22066 17816 22094
rect 17696 21729 17724 22066
rect 17682 21720 17738 21729
rect 17682 21655 17738 21664
rect 17696 16998 17724 21655
rect 17972 20466 18000 22374
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17880 19310 17908 20334
rect 18156 20058 18184 20742
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 18156 19446 18184 19722
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17866 17912 17922 17921
rect 17866 17847 17922 17856
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17696 15978 17724 16458
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17590 15056 17646 15065
rect 17590 14991 17646 15000
rect 17604 14958 17632 14991
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17696 14006 17724 15914
rect 17880 15502 17908 17847
rect 17972 16454 18000 18226
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 15162 18000 15302
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17868 14340 17920 14346
rect 18064 14328 18092 16934
rect 18156 14414 18184 19382
rect 18248 18358 18276 23530
rect 18340 21865 18368 24142
rect 18326 21856 18382 21865
rect 18326 21791 18382 21800
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18340 20754 18368 21422
rect 18432 20942 18460 25230
rect 18696 24608 18748 24614
rect 18696 24550 18748 24556
rect 18708 24274 18736 24550
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18708 23866 18736 24210
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18340 20726 18460 20754
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18340 19446 18368 19994
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18432 19334 18460 20726
rect 18340 19306 18460 19334
rect 18236 18352 18288 18358
rect 18236 18294 18288 18300
rect 18340 18170 18368 19306
rect 18524 18850 18552 23054
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18616 21350 18644 21490
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18604 19848 18656 19854
rect 18602 19816 18604 19825
rect 18656 19816 18658 19825
rect 18602 19751 18658 19760
rect 18432 18822 18552 18850
rect 18432 18698 18460 18822
rect 18420 18692 18472 18698
rect 18420 18634 18472 18640
rect 18248 18142 18368 18170
rect 18248 14618 18276 18142
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18340 16658 18368 18022
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18432 15502 18460 18634
rect 18800 17882 18828 23598
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18892 19446 18920 20198
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18524 15162 18552 15846
rect 18616 15366 18644 16526
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18708 15570 18736 15846
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18432 14822 18460 14962
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 17920 14300 18092 14328
rect 17868 14282 17920 14288
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17512 12434 17540 13806
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17512 12406 17632 12434
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17512 10470 17540 10678
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17420 9518 17448 9658
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17604 8922 17632 12406
rect 17420 8894 17632 8922
rect 17314 8664 17370 8673
rect 17314 8599 17370 8608
rect 17130 8256 17186 8265
rect 17130 8191 17186 8200
rect 17144 6866 17172 8191
rect 17328 7342 17356 8599
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17328 6866 17356 7278
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 17316 6724 17368 6730
rect 17316 6666 17368 6672
rect 17144 5846 17172 6666
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17236 6118 17264 6326
rect 17328 6322 17356 6666
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17420 5642 17448 8894
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17512 8634 17540 8774
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17512 7954 17540 8570
rect 17604 8498 17632 8774
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17590 8392 17646 8401
rect 17590 8327 17646 8336
rect 17604 7954 17632 8327
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17500 7744 17552 7750
rect 17696 7698 17724 12718
rect 17788 9654 17816 14214
rect 18156 14113 18184 14350
rect 18142 14104 18198 14113
rect 18142 14039 18198 14048
rect 17958 13560 18014 13569
rect 18248 13530 18276 14554
rect 18616 14482 18644 15302
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 14006 18736 14214
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18800 13870 18828 17818
rect 18892 15978 18920 19382
rect 18984 16114 19012 25706
rect 19076 20330 19104 26454
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19248 25832 19300 25838
rect 19248 25774 19300 25780
rect 19352 25786 19380 26318
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19444 25906 19472 26182
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19260 25294 19288 25774
rect 19352 25758 19472 25786
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19352 24818 19380 25638
rect 19444 24868 19472 25758
rect 19996 25430 20024 29582
rect 19984 25424 20036 25430
rect 19984 25366 20036 25372
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19444 24840 19564 24868
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 23730 19288 24006
rect 19248 23724 19300 23730
rect 19248 23666 19300 23672
rect 19352 22982 19380 24074
rect 19444 23497 19472 24686
rect 19536 24206 19564 24840
rect 20088 24410 20116 37198
rect 22112 36922 22140 37216
rect 22376 37188 22428 37194
rect 22376 37130 22428 37136
rect 22100 36916 22152 36922
rect 22100 36858 22152 36864
rect 22388 36854 22416 37130
rect 22376 36848 22428 36854
rect 22376 36790 22428 36796
rect 23216 36786 23244 39200
rect 24504 37126 24532 39200
rect 25148 37262 25176 39200
rect 26436 37262 26464 39200
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 25136 37256 25188 37262
rect 25136 37198 25188 37204
rect 26424 37256 26476 37262
rect 26424 37198 26476 37204
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 20628 36712 20680 36718
rect 20628 36654 20680 36660
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20168 26308 20220 26314
rect 20168 26250 20220 26256
rect 20180 24818 20208 26250
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19800 23860 19852 23866
rect 19800 23802 19852 23808
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19430 23488 19486 23497
rect 19430 23423 19486 23432
rect 19536 23186 19564 23598
rect 19812 23526 19840 23802
rect 20180 23730 20208 24618
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 19168 21622 19196 21898
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19246 18456 19302 18465
rect 19246 18391 19302 18400
rect 19260 18222 19288 18391
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18984 14482 19012 16050
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 17958 13495 18014 13504
rect 18236 13524 18288 13530
rect 17972 13190 18000 13495
rect 18236 13466 18288 13472
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17972 11830 18000 12582
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18064 11393 18092 13398
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18156 12345 18184 12378
rect 18142 12336 18198 12345
rect 18142 12271 18198 12280
rect 18616 11898 18644 13262
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 12918 18736 13126
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18800 12782 18828 13262
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18050 11384 18106 11393
rect 17960 11348 18012 11354
rect 18050 11319 18106 11328
rect 17960 11290 18012 11296
rect 17972 9722 18000 11290
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17788 9450 17816 9590
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17776 8968 17828 8974
rect 17774 8936 17776 8945
rect 17828 8936 17830 8945
rect 18064 8906 18092 9454
rect 17774 8871 17830 8880
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18156 8809 18184 8842
rect 18142 8800 18198 8809
rect 18142 8735 18198 8744
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17500 7686 17552 7692
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17420 5409 17448 5578
rect 17406 5400 17462 5409
rect 17406 5335 17462 5344
rect 17224 5160 17276 5166
rect 17052 5086 17172 5114
rect 17224 5102 17276 5108
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16776 3534 16804 3946
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16868 3482 16896 4218
rect 16960 3602 16988 4626
rect 17144 4434 17172 5086
rect 17052 4406 17172 4434
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 17052 3534 17080 4406
rect 17040 3528 17092 3534
rect 16776 3058 16804 3470
rect 16868 3454 16988 3482
rect 17040 3470 17092 3476
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16500 2876 16712 2904
rect 16500 2650 16528 2876
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16960 2446 16988 3454
rect 17236 2689 17264 5102
rect 17406 4992 17462 5001
rect 17406 4927 17462 4936
rect 17314 4856 17370 4865
rect 17314 4791 17370 4800
rect 17328 4486 17356 4791
rect 17420 4690 17448 4927
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 17222 2680 17278 2689
rect 17222 2615 17278 2624
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 15396 1834 15424 2382
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15488 2038 15516 2246
rect 15476 2032 15528 2038
rect 15476 1974 15528 1980
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 17328 1698 17356 2858
rect 17512 2650 17540 7686
rect 17604 7670 17724 7698
rect 17604 6730 17632 7670
rect 17682 7576 17738 7585
rect 17682 7511 17738 7520
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17590 6624 17646 6633
rect 17590 6559 17646 6568
rect 17604 6458 17632 6559
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17604 5273 17632 5306
rect 17590 5264 17646 5273
rect 17590 5199 17646 5208
rect 17696 5148 17724 7511
rect 17788 7342 17816 7890
rect 17880 7818 17908 8570
rect 18052 8560 18104 8566
rect 18104 8520 18184 8548
rect 18052 8502 18104 8508
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17960 7744 18012 7750
rect 17958 7712 17960 7721
rect 18012 7712 18014 7721
rect 17958 7647 18014 7656
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17604 5120 17724 5148
rect 17604 4078 17632 5120
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 17788 5001 17816 5034
rect 17774 4992 17830 5001
rect 17774 4927 17830 4936
rect 17682 4856 17738 4865
rect 17682 4791 17684 4800
rect 17736 4791 17738 4800
rect 17684 4762 17736 4768
rect 17682 4176 17738 4185
rect 17682 4111 17738 4120
rect 17696 4078 17724 4111
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17682 3904 17738 3913
rect 17682 3839 17738 3848
rect 17696 3398 17724 3839
rect 17788 3466 17816 4927
rect 17972 4690 18000 5714
rect 18064 4690 18092 8026
rect 18156 4826 18184 8520
rect 18248 8430 18276 10202
rect 18432 10062 18460 11086
rect 18694 10976 18750 10985
rect 18694 10911 18750 10920
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18524 10606 18552 10678
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18708 10130 18736 10911
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18892 10606 18920 10746
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18248 6730 18276 8026
rect 18432 8022 18460 9998
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18616 9674 18644 9930
rect 18984 9897 19012 12718
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19076 10198 19104 10542
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18970 9888 19026 9897
rect 18970 9823 19026 9832
rect 18616 9646 18736 9674
rect 18708 9178 18736 9646
rect 19168 9586 19196 9998
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18892 9110 18920 9386
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18524 8514 18552 9046
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18708 8673 18736 8910
rect 18694 8664 18750 8673
rect 18694 8599 18750 8608
rect 18616 8566 18644 8597
rect 18604 8560 18656 8566
rect 18524 8508 18604 8514
rect 18524 8502 18656 8508
rect 18524 8486 18644 8502
rect 18616 8430 18644 8486
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18340 7546 18368 7822
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 18248 2990 18276 6258
rect 18340 6254 18368 7278
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18340 5710 18368 6190
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18326 4312 18382 4321
rect 18326 4247 18382 4256
rect 18340 3058 18368 4247
rect 18432 3194 18460 7414
rect 18524 7206 18552 8366
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18524 6730 18552 7142
rect 18708 6769 18736 7142
rect 18694 6760 18750 6769
rect 18512 6724 18564 6730
rect 18694 6695 18750 6704
rect 18512 6666 18564 6672
rect 18510 6624 18566 6633
rect 18510 6559 18566 6568
rect 18524 6322 18552 6559
rect 18800 6390 18828 8978
rect 18880 8832 18932 8838
rect 18878 8800 18880 8809
rect 18932 8800 18934 8809
rect 18878 8735 18934 8744
rect 18984 8650 19012 9114
rect 18892 8622 19012 8650
rect 19062 8664 19118 8673
rect 18892 6730 18920 8622
rect 19062 8599 19118 8608
rect 19076 8430 19104 8599
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19156 7336 19208 7342
rect 19260 7324 19288 18158
rect 19352 16794 19380 19314
rect 19444 18970 19472 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21622 20024 23462
rect 20168 23044 20220 23050
rect 20168 22986 20220 22992
rect 20180 22166 20208 22986
rect 20272 22234 20300 31894
rect 20352 31136 20404 31142
rect 20352 31078 20404 31084
rect 20364 23662 20392 31078
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20168 22160 20220 22166
rect 20168 22102 20220 22108
rect 20352 22160 20404 22166
rect 20352 22102 20404 22108
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19800 21480 19852 21486
rect 19798 21448 19800 21457
rect 19852 21448 19854 21457
rect 20364 21418 20392 22102
rect 19798 21383 19854 21392
rect 20352 21412 20404 21418
rect 20352 21354 20404 21360
rect 20166 20904 20222 20913
rect 20166 20839 20222 20848
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19536 19854 19564 20266
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18154 20024 18702
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19444 16046 19472 17138
rect 19996 16590 20024 18090
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 14958 19380 15370
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19444 12730 19472 15982
rect 19996 15434 20024 16390
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19720 13734 19748 13806
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19720 13326 19748 13670
rect 20088 13530 20116 17546
rect 20180 17241 20208 20839
rect 20364 19786 20392 21354
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20272 18766 20300 19382
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 17746 20392 18566
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20166 17232 20222 17241
rect 20166 17167 20222 17176
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 15026 20208 16934
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20272 14482 20300 16390
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20364 14346 20392 15370
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20456 13852 20484 25978
rect 20536 21956 20588 21962
rect 20536 21898 20588 21904
rect 20548 21146 20576 21898
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20640 19446 20668 36654
rect 22284 35216 22336 35222
rect 22284 35158 22336 35164
rect 21364 34536 21416 34542
rect 21364 34478 21416 34484
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20548 14226 20576 18566
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20640 14618 20668 18294
rect 20732 15162 20760 28426
rect 20904 24676 20956 24682
rect 20904 24618 20956 24624
rect 20916 24342 20944 24618
rect 20904 24336 20956 24342
rect 20904 24278 20956 24284
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20824 16250 20852 16526
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20548 14198 20760 14226
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20180 13824 20484 13852
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20180 13410 20208 13824
rect 20548 13530 20576 14010
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20088 13382 20208 13410
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19616 12776 19668 12782
rect 19352 12702 19472 12730
rect 19614 12744 19616 12753
rect 19668 12744 19670 12753
rect 19352 11014 19380 12702
rect 19614 12679 19670 12688
rect 19628 12084 19656 12679
rect 19996 12646 20024 12922
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19444 12056 19656 12084
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19444 10742 19472 12056
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11121 20024 12106
rect 19982 11112 20038 11121
rect 19982 11047 20038 11056
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19982 10840 20038 10849
rect 19982 10775 20038 10784
rect 19432 10736 19484 10742
rect 19338 10704 19394 10713
rect 19996 10724 20024 10775
rect 19432 10678 19484 10684
rect 19904 10696 20024 10724
rect 19338 10639 19394 10648
rect 19352 8945 19380 10639
rect 19706 10432 19762 10441
rect 19706 10367 19762 10376
rect 19720 10266 19748 10367
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19444 9704 19472 10134
rect 19904 10130 19932 10696
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19996 10130 20024 10542
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19524 9988 19576 9994
rect 19892 9988 19944 9994
rect 19576 9948 19892 9976
rect 19524 9930 19576 9936
rect 19892 9930 19944 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19982 9752 20038 9761
rect 19444 9696 19982 9704
rect 19444 9687 20038 9696
rect 19444 9676 20024 9687
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19904 9382 19932 9454
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19996 9042 20024 9114
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19338 8936 19394 8945
rect 19338 8871 19394 8880
rect 19340 8832 19392 8838
rect 19338 8800 19340 8809
rect 19392 8800 19394 8809
rect 19338 8735 19394 8744
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19982 8664 20038 8673
rect 19708 8628 19760 8634
rect 19982 8599 20038 8608
rect 19708 8570 19760 8576
rect 19720 8514 19748 8570
rect 19996 8514 20024 8599
rect 20088 8548 20116 13382
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20180 8809 20208 13262
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20272 12434 20300 13194
rect 20364 12714 20392 13194
rect 20456 12714 20484 13398
rect 20732 13274 20760 14198
rect 20824 13938 20852 15574
rect 20916 15094 20944 16934
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20916 14550 20944 15030
rect 20904 14544 20956 14550
rect 20904 14486 20956 14492
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20916 13394 20944 14214
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20548 13246 20760 13274
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20352 12708 20404 12714
rect 20352 12650 20404 12656
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20272 12406 20392 12434
rect 20258 10432 20314 10441
rect 20258 10367 20314 10376
rect 20272 10198 20300 10367
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 20364 9874 20392 12406
rect 20548 12374 20576 13246
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12850 20760 13126
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20456 11694 20484 12106
rect 20640 11830 20668 12582
rect 20824 12102 20852 13262
rect 21008 13190 21036 13738
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 20996 12640 21048 12646
rect 21100 12617 21128 13738
rect 20996 12582 21048 12588
rect 21086 12608 21142 12617
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20272 9846 20392 9874
rect 20166 8800 20222 8809
rect 20166 8735 20222 8744
rect 20088 8520 20208 8548
rect 19720 8486 20024 8514
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19812 7954 19840 8366
rect 20076 8016 20128 8022
rect 20180 8004 20208 8520
rect 20272 8401 20300 9846
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20364 8974 20392 9658
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20352 8424 20404 8430
rect 20258 8392 20314 8401
rect 20352 8366 20404 8372
rect 20258 8327 20314 8336
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20128 7976 20208 8004
rect 20076 7958 20128 7964
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 20076 7880 20128 7886
rect 19890 7848 19946 7857
rect 20074 7848 20076 7857
rect 20168 7880 20220 7886
rect 20128 7848 20130 7857
rect 19946 7806 20024 7834
rect 19890 7783 19946 7792
rect 19996 7721 20024 7806
rect 20272 7868 20300 8026
rect 20364 7954 20392 8366
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20220 7840 20300 7868
rect 20168 7822 20220 7828
rect 20074 7783 20130 7792
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 20168 7744 20220 7750
rect 19982 7712 20038 7721
rect 20168 7686 20220 7692
rect 19574 7644 19882 7653
rect 19982 7647 20038 7656
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 19720 7342 19748 7414
rect 19208 7296 19288 7324
rect 19708 7336 19760 7342
rect 19156 7278 19208 7284
rect 19708 7278 19760 7284
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18616 6236 18644 6326
rect 18892 6236 18920 6666
rect 18616 6208 18920 6236
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18604 6112 18656 6118
rect 18984 6100 19012 6190
rect 18656 6072 19012 6100
rect 18604 6054 18656 6060
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18524 5642 18552 5714
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18524 3194 18552 5238
rect 18616 4622 18644 5782
rect 18696 5704 18748 5710
rect 18694 5672 18696 5681
rect 18748 5672 18750 5681
rect 18694 5607 18750 5616
rect 19076 5302 19104 7210
rect 19812 6916 19840 7278
rect 19352 6888 19840 6916
rect 19352 6882 19380 6888
rect 19168 6866 19380 6882
rect 19156 6860 19380 6866
rect 19208 6854 19380 6860
rect 19892 6860 19944 6866
rect 19156 6802 19208 6808
rect 19892 6802 19944 6808
rect 19340 6792 19392 6798
rect 19338 6760 19340 6769
rect 19392 6760 19394 6769
rect 19904 6746 19932 6802
rect 19720 6730 19932 6746
rect 19338 6695 19394 6704
rect 19708 6724 19932 6730
rect 19760 6718 19932 6724
rect 19708 6666 19760 6672
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19982 6624 20038 6633
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19168 5545 19196 6054
rect 19154 5536 19210 5545
rect 19154 5471 19210 5480
rect 19246 5400 19302 5409
rect 19246 5335 19302 5344
rect 18696 5296 18748 5302
rect 18696 5238 18748 5244
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 19156 5296 19208 5302
rect 19156 5238 19208 5244
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18708 3534 18736 5238
rect 18880 5092 18932 5098
rect 18880 5034 18932 5040
rect 18892 4826 18920 5034
rect 19168 5001 19196 5238
rect 19154 4992 19210 5001
rect 19154 4927 19210 4936
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 19156 4208 19208 4214
rect 19156 4150 19208 4156
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18984 3058 19012 3606
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 19076 2825 19104 4014
rect 19168 3194 19196 4150
rect 19260 4026 19288 5335
rect 19352 4978 19380 6598
rect 19574 6556 19882 6565
rect 19982 6559 20038 6568
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19800 6384 19852 6390
rect 19996 6372 20024 6559
rect 19852 6344 20024 6372
rect 19800 6326 19852 6332
rect 19432 5840 19484 5846
rect 19432 5782 19484 5788
rect 19444 5166 19472 5782
rect 19524 5704 19576 5710
rect 19522 5672 19524 5681
rect 19576 5672 19578 5681
rect 19522 5607 19578 5616
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20180 5409 20208 7686
rect 20364 7449 20392 7754
rect 20456 7721 20484 11222
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20536 11008 20588 11014
rect 20536 10950 20588 10956
rect 20548 9926 20576 10950
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20548 8362 20576 9454
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20442 7712 20498 7721
rect 20442 7647 20498 7656
rect 20548 7562 20576 8298
rect 20456 7534 20576 7562
rect 20456 7478 20484 7534
rect 20640 7478 20668 11018
rect 20732 9178 20760 11766
rect 20812 10736 20864 10742
rect 20916 10724 20944 12242
rect 21008 11082 21036 12582
rect 21086 12543 21142 12552
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 21100 11082 21128 12038
rect 21192 11626 21220 18362
rect 21284 17746 21312 19110
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 21270 15464 21326 15473
rect 21270 15399 21326 15408
rect 21284 15366 21312 15399
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 14618 21312 14962
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21284 12170 21312 12378
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21180 11620 21232 11626
rect 21180 11562 21232 11568
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21192 10742 21220 11562
rect 20864 10696 20944 10724
rect 21180 10736 21232 10742
rect 20812 10678 20864 10684
rect 21180 10678 21232 10684
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20996 10464 21048 10470
rect 20994 10432 20996 10441
rect 21048 10432 21050 10441
rect 20994 10367 21050 10376
rect 21100 9722 21128 10542
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20732 8090 20760 8434
rect 20824 8090 20852 8842
rect 20916 8430 20944 8978
rect 21192 8906 21220 10406
rect 21284 10033 21312 10678
rect 21270 10024 21326 10033
rect 21270 9959 21326 9968
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21008 8430 21036 8570
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20444 7472 20496 7478
rect 20350 7440 20406 7449
rect 20444 7414 20496 7420
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20350 7375 20406 7384
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20272 6798 20300 7278
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20732 6458 20760 7890
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20352 6112 20404 6118
rect 20352 6054 20404 6060
rect 20260 5840 20312 5846
rect 20260 5782 20312 5788
rect 20166 5400 20222 5409
rect 20166 5335 20222 5344
rect 19708 5296 19760 5302
rect 19760 5256 20024 5284
rect 19708 5238 19760 5244
rect 19996 5166 20024 5256
rect 19432 5160 19484 5166
rect 19892 5160 19944 5166
rect 19484 5108 19564 5114
rect 19432 5102 19564 5108
rect 19892 5102 19944 5108
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19444 5086 19564 5102
rect 19430 4992 19486 5001
rect 19352 4950 19430 4978
rect 19430 4927 19486 4936
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19352 4185 19380 4694
rect 19444 4690 19472 4927
rect 19536 4826 19564 5086
rect 19904 5030 19932 5102
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19536 4536 19564 4762
rect 19444 4508 19564 4536
rect 19444 4282 19472 4508
rect 19904 4486 19932 4762
rect 20168 4684 20220 4690
rect 20272 4672 20300 5782
rect 20364 5710 20392 6054
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20442 5536 20498 5545
rect 20442 5471 20498 5480
rect 20456 5234 20484 5471
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20548 4826 20576 6326
rect 20640 6254 20668 6394
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20640 5114 20668 5306
rect 20732 5234 20760 5850
rect 20824 5302 20852 7890
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20916 5778 20944 7482
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20902 5400 20958 5409
rect 20902 5335 20958 5344
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20812 5160 20864 5166
rect 20640 5086 20760 5114
rect 20812 5102 20864 5108
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20364 4706 20392 4762
rect 20364 4678 20484 4706
rect 20220 4644 20300 4672
rect 20168 4626 20220 4632
rect 20352 4616 20404 4622
rect 20456 4593 20484 4678
rect 20352 4558 20404 4564
rect 20442 4584 20498 4593
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19338 4176 19394 4185
rect 19996 4146 20024 4422
rect 20166 4312 20222 4321
rect 20364 4282 20392 4558
rect 20442 4519 20498 4528
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20166 4247 20222 4256
rect 20352 4276 20404 4282
rect 19338 4111 19394 4120
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19260 3998 19380 4026
rect 19352 3602 19380 3998
rect 20180 3738 20208 4247
rect 20352 4218 20404 4224
rect 20548 4146 20576 4490
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20534 4040 20590 4049
rect 20534 3975 20590 3984
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19904 3482 19932 3674
rect 20076 3664 20128 3670
rect 20352 3664 20404 3670
rect 20128 3612 20352 3618
rect 20076 3606 20404 3612
rect 20088 3590 20392 3606
rect 20548 3602 20576 3975
rect 20640 3738 20668 4966
rect 20732 4282 20760 5086
rect 20720 4276 20772 4282
rect 20720 4218 20772 4224
rect 20718 4176 20774 4185
rect 20718 4111 20774 4120
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19062 2816 19118 2825
rect 19062 2751 19118 2760
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17972 2038 18000 2314
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 17960 2032 18012 2038
rect 17960 1974 18012 1980
rect 16120 1692 16172 1698
rect 16120 1634 16172 1640
rect 17316 1692 17368 1698
rect 17316 1634 17368 1640
rect 17408 1692 17460 1698
rect 17408 1634 17460 1640
rect 14832 1284 14884 1290
rect 14832 1226 14884 1232
rect 14844 800 14872 1226
rect 16132 800 16160 1634
rect 17420 800 17448 1634
rect 18064 800 18092 2246
rect 19260 1902 19288 2450
rect 19248 1896 19300 1902
rect 19248 1838 19300 1844
rect 19352 800 19380 2926
rect 19444 2582 19472 3470
rect 19708 3460 19760 3466
rect 19904 3454 20392 3482
rect 19760 3420 19840 3448
rect 19708 3402 19760 3408
rect 19812 3380 19840 3420
rect 20076 3392 20128 3398
rect 19812 3352 20024 3380
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3097 20024 3352
rect 20074 3360 20076 3369
rect 20128 3360 20130 3369
rect 20074 3295 20130 3304
rect 20166 3224 20222 3233
rect 20166 3159 20222 3168
rect 19614 3088 19670 3097
rect 19614 3023 19616 3032
rect 19668 3023 19670 3032
rect 19982 3088 20038 3097
rect 20180 3058 20208 3159
rect 20364 3058 20392 3454
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 20548 3369 20576 3402
rect 20732 3369 20760 4111
rect 20824 4010 20852 5102
rect 20916 4321 20944 5335
rect 20902 4312 20958 4321
rect 20902 4247 20958 4256
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20534 3360 20590 3369
rect 20534 3295 20590 3304
rect 20718 3360 20774 3369
rect 20718 3295 20774 3304
rect 20824 3194 20852 3538
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 19982 3023 20038 3032
rect 20168 3052 20220 3058
rect 19616 2994 19668 3000
rect 20168 2994 20220 3000
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20180 2961 20208 2994
rect 20166 2952 20222 2961
rect 20166 2887 20222 2896
rect 20350 2952 20406 2961
rect 20350 2887 20406 2896
rect 20536 2916 20588 2922
rect 20364 2650 20392 2887
rect 20536 2858 20588 2864
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20088 1970 20116 2382
rect 20076 1964 20128 1970
rect 20076 1906 20128 1912
rect 20548 1358 20576 2858
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20536 1352 20588 1358
rect 20536 1294 20588 1300
rect 20640 800 20668 2382
rect 21008 2310 21036 7414
rect 21100 6322 21128 8434
rect 21192 7954 21220 8842
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21284 7478 21312 9590
rect 21376 8566 21404 34478
rect 21916 25152 21968 25158
rect 21916 25094 21968 25100
rect 21928 24750 21956 25094
rect 22192 24880 22244 24886
rect 22192 24822 22244 24828
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 22204 24614 22232 24822
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 21468 19514 21496 19722
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 16522 21496 17478
rect 21456 16516 21508 16522
rect 21456 16458 21508 16464
rect 21468 14550 21496 16458
rect 21560 15638 21588 22578
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21744 21554 21772 21830
rect 22204 21554 22232 22918
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21640 19984 21692 19990
rect 21640 19926 21692 19932
rect 21652 19786 21680 19926
rect 21640 19780 21692 19786
rect 21640 19722 21692 19728
rect 21744 16674 21772 20946
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 21928 18222 21956 19178
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21652 16646 21772 16674
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21560 15366 21588 15574
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 12434 21588 14350
rect 21468 12406 21588 12434
rect 21468 9024 21496 12406
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21560 11762 21588 12106
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21652 11558 21680 16646
rect 21824 16040 21876 16046
rect 21824 15982 21876 15988
rect 21732 15972 21784 15978
rect 21732 15914 21784 15920
rect 21744 15706 21772 15914
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 21744 12102 21772 15642
rect 21836 15502 21864 15982
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15094 21864 15438
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21928 14414 21956 18158
rect 22204 16590 22232 19314
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22020 15348 22048 16390
rect 22192 16176 22244 16182
rect 22192 16118 22244 16124
rect 22020 15320 22140 15348
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 14482 22048 14962
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 22112 13870 22140 15320
rect 22204 15162 22232 16118
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21744 11354 21772 11494
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21836 11268 21864 12786
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21928 11608 21956 12174
rect 22112 11898 22140 12582
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 21928 11580 22048 11608
rect 21916 11280 21968 11286
rect 21836 11240 21916 11268
rect 21916 11222 21968 11228
rect 21914 11112 21970 11121
rect 21914 11047 21916 11056
rect 21968 11047 21970 11056
rect 21916 11018 21968 11024
rect 22020 10742 22048 11580
rect 22204 11218 22232 11630
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22008 10736 22060 10742
rect 21546 10704 21602 10713
rect 22008 10678 22060 10684
rect 21546 10639 21548 10648
rect 21600 10639 21602 10648
rect 21548 10610 21600 10616
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22112 10441 22140 10542
rect 22098 10432 22154 10441
rect 22098 10367 22154 10376
rect 22296 10266 22324 35158
rect 24596 34542 24624 37198
rect 27724 37126 27752 39200
rect 28368 37262 28396 39200
rect 29656 37262 29684 39200
rect 30944 37330 30972 39200
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 24584 34536 24636 34542
rect 24584 34478 24636 34484
rect 25332 31890 25360 37062
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 25320 31884 25372 31890
rect 25320 31826 25372 31832
rect 26252 31346 26280 36722
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22848 25362 22876 26182
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22848 24206 22876 24754
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23308 23118 23336 23462
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23492 22642 23520 23666
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22388 20874 22416 21286
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22388 20602 22416 20810
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22572 20330 22600 21830
rect 23124 21486 23152 22034
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23112 21480 23164 21486
rect 23112 21422 23164 21428
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22480 14074 22508 15642
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21652 9466 21680 10066
rect 21822 10024 21878 10033
rect 21822 9959 21824 9968
rect 21876 9959 21878 9968
rect 22100 9988 22152 9994
rect 21824 9930 21876 9936
rect 22100 9930 22152 9936
rect 22112 9674 22140 9930
rect 22020 9646 22140 9674
rect 22388 9654 22416 13874
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22480 13530 22508 13806
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22572 12646 22600 20266
rect 23400 19922 23428 21490
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23676 20602 23704 21422
rect 23756 21072 23808 21078
rect 23756 21014 23808 21020
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22848 18698 22876 18906
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22480 11558 22508 12038
rect 22572 11665 22600 12174
rect 22558 11656 22614 11665
rect 22558 11591 22614 11600
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22572 10674 22600 11494
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22664 10554 22692 17750
rect 22848 13394 22876 18634
rect 23216 18426 23244 18634
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23400 18290 23428 19110
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23584 18222 23612 20402
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23768 17202 23796 21014
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 23860 20602 23888 20810
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 24044 19922 24072 28018
rect 24872 26450 24900 28358
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24124 25288 24176 25294
rect 24124 25230 24176 25236
rect 24136 21078 24164 25230
rect 26252 24682 26280 27406
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23952 19514 23980 19654
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24044 18834 24072 19858
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23846 17096 23902 17105
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22940 15434 22968 16526
rect 23032 15706 23060 17070
rect 23846 17031 23902 17040
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23400 15638 23428 16458
rect 23388 15632 23440 15638
rect 23388 15574 23440 15580
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 23860 15026 23888 17031
rect 23952 16590 23980 17206
rect 24044 17066 24072 18226
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24044 16658 24072 17002
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23202 14512 23258 14521
rect 23202 14447 23258 14456
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22756 12918 22784 13194
rect 22744 12912 22796 12918
rect 22744 12854 22796 12860
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22848 11082 22876 12582
rect 22940 12434 22968 13670
rect 22940 12406 23060 12434
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22572 10526 22692 10554
rect 22376 9648 22428 9654
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21652 9438 21772 9466
rect 21468 8996 21588 9024
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21468 8566 21496 8842
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21456 8560 21508 8566
rect 21456 8502 21508 8508
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21192 6458 21220 6598
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21284 6066 21312 7278
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21100 6038 21312 6066
rect 21100 5710 21128 6038
rect 21270 5944 21326 5953
rect 21270 5879 21326 5888
rect 21178 5808 21234 5817
rect 21178 5743 21234 5752
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 21088 5296 21140 5302
rect 21088 5238 21140 5244
rect 21192 5250 21220 5743
rect 21284 5409 21312 5879
rect 21376 5817 21404 6666
rect 21456 6384 21508 6390
rect 21456 6326 21508 6332
rect 21362 5808 21418 5817
rect 21362 5743 21418 5752
rect 21468 5574 21496 6326
rect 21560 5710 21588 8996
rect 21744 8906 21772 9438
rect 21732 8900 21784 8906
rect 21732 8842 21784 8848
rect 21730 8392 21786 8401
rect 21730 8327 21786 8336
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21652 7546 21680 7754
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21652 5914 21680 6870
rect 21744 6322 21772 8327
rect 21836 7954 21864 9522
rect 21928 8838 21956 9522
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 22020 8537 22048 9646
rect 22376 9590 22428 9596
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22112 8634 22140 9318
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22006 8528 22062 8537
rect 22006 8463 22008 8472
rect 22060 8463 22062 8472
rect 22008 8434 22060 8440
rect 22388 8362 22416 9590
rect 22572 9194 22600 10526
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22940 10266 22968 10406
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22756 9654 22784 9862
rect 22834 9752 22890 9761
rect 22834 9687 22890 9696
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22572 9166 22784 9194
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22466 8120 22522 8129
rect 22466 8055 22522 8064
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 22374 7848 22430 7857
rect 21824 7812 21876 7818
rect 22374 7783 22430 7792
rect 21824 7754 21876 7760
rect 21836 7274 21864 7754
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 22020 7041 22048 7346
rect 22006 7032 22062 7041
rect 22006 6967 22062 6976
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 22008 6656 22060 6662
rect 22192 6656 22244 6662
rect 22060 6616 22192 6644
rect 22008 6598 22060 6604
rect 22192 6598 22244 6604
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21744 5710 21772 6258
rect 21836 6186 21864 6598
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21822 6080 21878 6089
rect 21822 6015 21878 6024
rect 21548 5704 21600 5710
rect 21732 5704 21784 5710
rect 21548 5646 21600 5652
rect 21638 5672 21694 5681
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21270 5400 21326 5409
rect 21270 5335 21326 5344
rect 21100 5137 21128 5238
rect 21192 5234 21312 5250
rect 21192 5228 21324 5234
rect 21192 5222 21272 5228
rect 21272 5170 21324 5176
rect 21086 5128 21142 5137
rect 21086 5063 21142 5072
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 21100 3466 21128 4490
rect 21192 4078 21220 4966
rect 21284 4690 21312 4966
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21376 4486 21404 4762
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 21284 1222 21312 4014
rect 21468 3534 21496 5510
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21376 3194 21404 3470
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21560 1630 21588 5646
rect 21836 5681 21864 6015
rect 21732 5646 21784 5652
rect 21822 5672 21878 5681
rect 21638 5607 21694 5616
rect 21822 5607 21878 5616
rect 21652 4486 21680 5607
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21730 5400 21786 5409
rect 21730 5335 21786 5344
rect 21640 4480 21692 4486
rect 21640 4422 21692 4428
rect 21744 4010 21772 5335
rect 21732 4004 21784 4010
rect 21732 3946 21784 3952
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21652 2825 21680 3878
rect 21836 3641 21864 5510
rect 21822 3632 21878 3641
rect 21928 3602 21956 6326
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 5001 22048 6054
rect 22112 5545 22140 6258
rect 22388 5658 22416 7783
rect 22480 6610 22508 8055
rect 22572 7750 22600 8774
rect 22664 7886 22692 9046
rect 22756 8974 22784 9166
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22480 6582 22600 6610
rect 22572 6458 22600 6582
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22480 5710 22508 6394
rect 22204 5630 22416 5658
rect 22468 5704 22520 5710
rect 22468 5646 22520 5652
rect 22098 5536 22154 5545
rect 22098 5471 22154 5480
rect 22006 4992 22062 5001
rect 22006 4927 22062 4936
rect 22008 4752 22060 4758
rect 22006 4720 22008 4729
rect 22060 4720 22062 4729
rect 22006 4655 22062 4664
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 4282 22048 4422
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22204 4146 22232 5630
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22100 3664 22152 3670
rect 22098 3632 22100 3641
rect 22152 3632 22154 3641
rect 21822 3567 21878 3576
rect 21916 3596 21968 3602
rect 22098 3567 22154 3576
rect 21916 3538 21968 3544
rect 22192 3392 22244 3398
rect 22112 3352 22192 3380
rect 21914 2952 21970 2961
rect 21914 2887 21970 2896
rect 21928 2854 21956 2887
rect 21824 2848 21876 2854
rect 21638 2816 21694 2825
rect 21824 2790 21876 2796
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21638 2751 21694 2760
rect 21836 2514 21864 2790
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 21548 1624 21600 1630
rect 21548 1566 21600 1572
rect 21272 1216 21324 1222
rect 21272 1158 21324 1164
rect 21928 800 21956 2382
rect 22112 1873 22140 3352
rect 22192 3334 22244 3340
rect 22296 3210 22324 5238
rect 22204 3182 22324 3210
rect 22098 1864 22154 1873
rect 22098 1799 22154 1808
rect 22204 1766 22232 3182
rect 22388 3126 22416 5510
rect 22664 5386 22692 6734
rect 22572 5358 22692 5386
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22480 4622 22508 5170
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22376 3120 22428 3126
rect 22480 3097 22508 3470
rect 22376 3062 22428 3068
rect 22466 3088 22522 3097
rect 22466 3023 22522 3032
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22296 1766 22324 2926
rect 22572 2825 22600 5358
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22664 3233 22692 5170
rect 22756 5137 22784 8910
rect 22848 6254 22876 9687
rect 23032 7546 23060 12406
rect 23216 12238 23244 14447
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 23308 12850 23336 13738
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23400 13326 23428 13670
rect 23388 13320 23440 13326
rect 23584 13297 23612 13874
rect 23940 13320 23992 13326
rect 23388 13262 23440 13268
rect 23570 13288 23626 13297
rect 23940 13262 23992 13268
rect 23570 13223 23626 13232
rect 23388 12912 23440 12918
rect 23386 12880 23388 12889
rect 23440 12880 23442 12889
rect 23296 12844 23348 12850
rect 23386 12815 23442 12824
rect 23296 12786 23348 12792
rect 23294 12472 23350 12481
rect 23294 12407 23296 12416
rect 23348 12407 23350 12416
rect 23296 12378 23348 12384
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23112 11824 23164 11830
rect 23112 11766 23164 11772
rect 23294 11792 23350 11801
rect 23124 11626 23152 11766
rect 23584 11762 23612 13223
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23676 12434 23704 13126
rect 23952 12986 23980 13262
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23676 12406 23796 12434
rect 23294 11727 23350 11736
rect 23572 11756 23624 11762
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23308 11150 23336 11727
rect 23572 11698 23624 11704
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 23124 10538 23152 11018
rect 23294 10568 23350 10577
rect 23112 10532 23164 10538
rect 23294 10503 23350 10512
rect 23112 10474 23164 10480
rect 23124 9586 23152 10474
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23204 9444 23256 9450
rect 23204 9386 23256 9392
rect 23110 9208 23166 9217
rect 23110 9143 23166 9152
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22926 7440 22982 7449
rect 22926 7375 22982 7384
rect 22940 6322 22968 7375
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22742 5128 22798 5137
rect 22742 5063 22798 5072
rect 22836 5024 22888 5030
rect 22836 4966 22888 4972
rect 22742 4312 22798 4321
rect 22742 4247 22744 4256
rect 22796 4247 22798 4256
rect 22744 4218 22796 4224
rect 22848 3913 22876 4966
rect 22834 3904 22890 3913
rect 22834 3839 22890 3848
rect 22650 3224 22706 3233
rect 22650 3159 22706 3168
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22558 2816 22614 2825
rect 22558 2751 22614 2760
rect 22664 2650 22692 2994
rect 22940 2990 22968 6258
rect 23124 5710 23152 9143
rect 23216 7886 23244 9386
rect 23308 8378 23336 10503
rect 23662 10296 23718 10305
rect 23662 10231 23718 10240
rect 23386 9344 23442 9353
rect 23386 9279 23442 9288
rect 23400 9042 23428 9279
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23400 8498 23428 8978
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23308 8350 23428 8378
rect 23400 7886 23428 8350
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23112 5704 23164 5710
rect 23032 5664 23112 5692
rect 23032 4078 23060 5664
rect 23112 5646 23164 5652
rect 23216 4826 23244 6938
rect 23400 6866 23428 7278
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23492 6798 23520 7142
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23584 6458 23612 6734
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23308 5681 23336 6258
rect 23570 6216 23626 6225
rect 23570 6151 23626 6160
rect 23294 5672 23350 5681
rect 23294 5607 23350 5616
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 23400 4865 23428 5170
rect 23480 5092 23532 5098
rect 23480 5034 23532 5040
rect 23386 4856 23442 4865
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23204 4820 23256 4826
rect 23386 4791 23442 4800
rect 23204 4762 23256 4768
rect 23124 4622 23152 4762
rect 23492 4706 23520 5034
rect 23400 4690 23520 4706
rect 23388 4684 23520 4690
rect 23440 4678 23520 4684
rect 23388 4626 23440 4632
rect 23584 4622 23612 6151
rect 23676 5846 23704 10231
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23112 4616 23164 4622
rect 23296 4616 23348 4622
rect 23164 4576 23244 4604
rect 23112 4558 23164 4564
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 23124 4282 23152 4422
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23216 4078 23244 4576
rect 23296 4558 23348 4564
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23662 4584 23718 4593
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23308 3777 23336 4558
rect 23662 4519 23664 4528
rect 23716 4519 23718 4528
rect 23664 4490 23716 4496
rect 23768 4146 23796 12406
rect 24032 11756 24084 11762
rect 24032 11698 24084 11704
rect 23846 10024 23902 10033
rect 23846 9959 23848 9968
rect 23900 9959 23902 9968
rect 23848 9930 23900 9936
rect 24044 9586 24072 11698
rect 24122 10840 24178 10849
rect 24122 10775 24124 10784
rect 24176 10775 24178 10784
rect 24124 10746 24176 10752
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24228 10130 24256 10542
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23846 9480 23902 9489
rect 23846 9415 23902 9424
rect 23860 9178 23888 9415
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23846 7576 23902 7585
rect 23846 7511 23902 7520
rect 23860 4622 23888 7511
rect 23952 6633 23980 8910
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 23938 6624 23994 6633
rect 23938 6559 23994 6568
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23294 3768 23350 3777
rect 23294 3703 23350 3712
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 22756 2689 22784 2790
rect 22742 2680 22798 2689
rect 22652 2644 22704 2650
rect 22742 2615 22798 2624
rect 22652 2586 22704 2592
rect 23308 2378 23336 2790
rect 23400 2553 23428 3878
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2582 23520 3334
rect 23480 2576 23532 2582
rect 23386 2544 23442 2553
rect 23480 2518 23532 2524
rect 23386 2479 23442 2488
rect 23572 2440 23624 2446
rect 23386 2408 23442 2417
rect 23296 2372 23348 2378
rect 23572 2382 23624 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 23386 2343 23442 2352
rect 23296 2314 23348 2320
rect 23400 2310 23428 2343
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 23388 2304 23440 2310
rect 23388 2246 23440 2252
rect 22192 1760 22244 1766
rect 22192 1702 22244 1708
rect 22284 1760 22336 1766
rect 22284 1702 22336 1708
rect 22572 800 22600 2246
rect 23584 1698 23612 2382
rect 23572 1692 23624 1698
rect 23572 1634 23624 1640
rect 23860 800 23888 2382
rect 23952 1737 23980 6258
rect 24044 5234 24072 7890
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 23938 1728 23994 1737
rect 23938 1663 23994 1672
rect 24044 1601 24072 3878
rect 24136 1902 24164 3878
rect 24228 3534 24256 7346
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 2990 24256 3470
rect 24216 2984 24268 2990
rect 24216 2926 24268 2932
rect 24320 2650 24348 24142
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24398 21448 24454 21457
rect 24398 21383 24454 21392
rect 24412 21350 24440 21383
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 24412 18426 24440 20402
rect 24596 19854 24624 23598
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 25424 21690 25452 21898
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 26240 21616 26292 21622
rect 26240 21558 26292 21564
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24872 20398 24900 20742
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24964 19446 24992 19654
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24412 16454 24440 17070
rect 24872 16658 24900 19246
rect 24964 18834 24992 19246
rect 25148 19145 25176 21490
rect 26252 21146 26280 21558
rect 26332 21412 26384 21418
rect 26332 21354 26384 21360
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26344 21146 26372 21354
rect 26240 21140 26292 21146
rect 26240 21082 26292 21088
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 25792 20058 25820 20470
rect 26528 20398 26556 21354
rect 26712 20602 26740 31078
rect 27172 30734 27200 37062
rect 27816 36922 27844 37198
rect 31300 37188 31352 37194
rect 31300 37130 31352 37136
rect 28540 37120 28592 37126
rect 28540 37062 28592 37068
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 28552 32910 28580 37062
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28644 31822 28672 37062
rect 31312 36786 31340 37130
rect 32232 37126 32260 39200
rect 32876 37262 32904 39200
rect 34164 37330 34192 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37346 35480 39200
rect 34152 37324 34204 37330
rect 35452 37318 35572 37346
rect 34152 37266 34204 37272
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32864 37256 32916 37262
rect 32864 37198 32916 37204
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 31300 36780 31352 36786
rect 31300 36722 31352 36728
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 27160 30728 27212 30734
rect 27160 30670 27212 30676
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31772 27606 31800 29106
rect 31760 27600 31812 27606
rect 31760 27542 31812 27548
rect 31116 25492 31168 25498
rect 31116 25434 31168 25440
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 29104 23866 29132 24550
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 29012 22098 29040 23462
rect 29736 22772 29788 22778
rect 29736 22714 29788 22720
rect 29000 22092 29052 22098
rect 29000 22034 29052 22040
rect 26792 20800 26844 20806
rect 26792 20742 26844 20748
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 25780 20052 25832 20058
rect 25780 19994 25832 20000
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 25516 19446 25544 19926
rect 26804 19854 26832 20742
rect 26976 20392 27028 20398
rect 26976 20334 27028 20340
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26896 19922 26924 20198
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26988 19854 27016 20334
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25134 19136 25190 19145
rect 25134 19071 25190 19080
rect 25686 19136 25742 19145
rect 25686 19071 25742 19080
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25056 18426 25084 18702
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 25700 18290 25728 19071
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25780 18080 25832 18086
rect 25780 18022 25832 18028
rect 25792 17270 25820 18022
rect 25780 17264 25832 17270
rect 25780 17206 25832 17212
rect 25688 17128 25740 17134
rect 25688 17070 25740 17076
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24780 16250 24808 16458
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24596 15570 24624 15982
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24780 15570 24808 15846
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24674 14648 24730 14657
rect 24674 14583 24730 14592
rect 24492 10464 24544 10470
rect 24492 10406 24544 10412
rect 24398 9616 24454 9625
rect 24504 9586 24532 10406
rect 24398 9551 24454 9560
rect 24492 9580 24544 9586
rect 24412 6390 24440 9551
rect 24492 9522 24544 9528
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24596 9178 24624 9522
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24688 6798 24716 14583
rect 24780 14482 24808 14758
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24858 12200 24914 12209
rect 24858 12135 24914 12144
rect 24872 11898 24900 12135
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24780 11354 24808 11698
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24780 10062 24808 10950
rect 25042 10160 25098 10169
rect 25042 10095 25098 10104
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24872 8362 24900 9318
rect 25056 8498 25084 10095
rect 25516 9178 25544 16594
rect 25700 16522 25728 17070
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 26160 16658 26188 16934
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 27712 16652 27764 16658
rect 27712 16594 27764 16600
rect 25688 16516 25740 16522
rect 25688 16458 25740 16464
rect 25700 15978 25728 16458
rect 26792 16448 26844 16454
rect 26792 16390 26844 16396
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 25688 15972 25740 15978
rect 25688 15914 25740 15920
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25884 10742 25912 13262
rect 25964 11008 26016 11014
rect 25964 10950 26016 10956
rect 25872 10736 25924 10742
rect 25872 10678 25924 10684
rect 25976 10674 26004 10950
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 26068 10062 26096 14962
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 26160 14414 26188 14894
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26252 13462 26280 16050
rect 26804 15706 26832 16390
rect 27724 16250 27752 16594
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27618 16144 27674 16153
rect 27618 16079 27620 16088
rect 27672 16079 27674 16088
rect 27620 16050 27672 16056
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 27988 15632 28040 15638
rect 27988 15574 28040 15580
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26712 14482 26740 14894
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26608 14272 26660 14278
rect 26608 14214 26660 14220
rect 26620 14074 26648 14214
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26620 13870 26648 14010
rect 26804 14006 26832 14758
rect 28000 14414 28028 15574
rect 28816 15360 28868 15366
rect 28816 15302 28868 15308
rect 28828 15026 28856 15302
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27344 14272 27396 14278
rect 27344 14214 27396 14220
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 26792 14000 26844 14006
rect 26792 13942 26844 13948
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26804 13530 26832 13942
rect 27356 13938 27384 14214
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 27252 13456 27304 13462
rect 27252 13398 27304 13404
rect 27264 13326 27292 13398
rect 28092 13394 28120 14214
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27344 13184 27396 13190
rect 27344 13126 27396 13132
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26160 11150 26188 11494
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 26148 11144 26200 11150
rect 26148 11086 26200 11092
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26620 10606 26648 10950
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25504 9172 25556 9178
rect 25504 9114 25556 9120
rect 25226 9072 25282 9081
rect 25226 9007 25282 9016
rect 25240 8974 25268 9007
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25332 8673 25360 8774
rect 25318 8664 25374 8673
rect 25318 8599 25374 8608
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24400 6384 24452 6390
rect 24688 6361 24716 6598
rect 24400 6326 24452 6332
rect 24674 6352 24730 6361
rect 24674 6287 24730 6296
rect 24780 4842 24808 8230
rect 25056 7410 25084 8434
rect 25226 7984 25282 7993
rect 25226 7919 25282 7928
rect 25240 7546 25268 7919
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 24860 7336 24912 7342
rect 24858 7304 24860 7313
rect 24912 7304 24914 7313
rect 24858 7239 24914 7248
rect 24858 7168 24914 7177
rect 24858 7103 24914 7112
rect 24872 5914 24900 7103
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 25056 5846 25084 7346
rect 25596 6112 25648 6118
rect 25596 6054 25648 6060
rect 25044 5840 25096 5846
rect 25044 5782 25096 5788
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 24492 4820 24544 4826
rect 24780 4814 24900 4842
rect 24492 4762 24544 4768
rect 24504 4622 24532 4762
rect 24872 4758 24900 4814
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 24780 4486 24808 4626
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24596 3534 24624 4422
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24596 2922 24624 3470
rect 24688 3126 24716 3674
rect 24676 3120 24728 3126
rect 24676 3062 24728 3068
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 24308 2644 24360 2650
rect 24308 2586 24360 2592
rect 24124 1896 24176 1902
rect 24124 1838 24176 1844
rect 24030 1592 24086 1601
rect 24030 1527 24086 1536
rect 24780 1290 24808 3946
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24872 2038 24900 3334
rect 24860 2032 24912 2038
rect 24860 1974 24912 1980
rect 24768 1284 24820 1290
rect 24768 1226 24820 1232
rect 12898 200 12954 800
rect 14186 200 14242 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 17406 200 17462 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 21914 200 21970 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 24964 202 24992 5170
rect 25412 5092 25464 5098
rect 25412 5034 25464 5040
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 25056 3602 25084 4422
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 25148 3534 25176 4014
rect 25136 3528 25188 3534
rect 25136 3470 25188 3476
rect 25424 3058 25452 5034
rect 25502 4448 25558 4457
rect 25502 4383 25558 4392
rect 25516 3126 25544 4383
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25332 2650 25360 2994
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 25608 2446 25636 6054
rect 25870 5264 25926 5273
rect 25870 5199 25926 5208
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25792 3534 25820 4082
rect 25884 3738 25912 5199
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25148 800 25176 2246
rect 25700 1358 25728 2994
rect 25976 2446 26004 9862
rect 26148 8356 26200 8362
rect 26148 8298 26200 8304
rect 26054 6896 26110 6905
rect 26054 6831 26110 6840
rect 26068 2854 26096 6831
rect 26160 6322 26188 8298
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 26436 5914 26464 6258
rect 26424 5908 26476 5914
rect 26424 5850 26476 5856
rect 26896 4010 26924 11222
rect 27356 11121 27384 13126
rect 27342 11112 27398 11121
rect 27342 11047 27398 11056
rect 28264 9988 28316 9994
rect 28264 9930 28316 9936
rect 28170 5808 28226 5817
rect 28170 5743 28226 5752
rect 28184 4826 28212 5743
rect 28276 4826 28304 9930
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 28172 4820 28224 4826
rect 28172 4762 28224 4768
rect 28264 4820 28316 4826
rect 28264 4762 28316 4768
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 26884 4004 26936 4010
rect 26884 3946 26936 3952
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26608 3392 26660 3398
rect 26606 3360 26608 3369
rect 26660 3360 26662 3369
rect 26606 3295 26662 3304
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25688 1352 25740 1358
rect 25688 1294 25740 1300
rect 25792 800 25820 2246
rect 26712 1970 26740 3878
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 26700 1964 26752 1970
rect 26700 1906 26752 1912
rect 27080 800 27108 2382
rect 27172 2009 27200 3334
rect 27252 2848 27304 2854
rect 27252 2790 27304 2796
rect 27264 2106 27292 2790
rect 27252 2100 27304 2106
rect 27252 2042 27304 2048
rect 27158 2000 27214 2009
rect 27158 1935 27214 1944
rect 24952 196 25004 202
rect 25134 200 25190 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 24952 138 25004 144
rect 11704 128 11756 134
rect 11704 70 11756 76
rect 27356 66 27384 4082
rect 27986 3632 28042 3641
rect 27986 3567 28042 3576
rect 28000 3534 28028 3567
rect 27988 3528 28040 3534
rect 27802 3496 27858 3505
rect 27436 3460 27488 3466
rect 27988 3470 28040 3476
rect 27802 3431 27858 3440
rect 27436 3402 27488 3408
rect 27448 2990 27476 3402
rect 27816 3398 27844 3431
rect 27804 3392 27856 3398
rect 27804 3334 27856 3340
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 27436 2984 27488 2990
rect 27436 2926 27488 2932
rect 28000 134 28028 2994
rect 28460 2650 28488 6190
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 29748 2446 29776 22714
rect 30472 21548 30524 21554
rect 30472 21490 30524 21496
rect 29920 21004 29972 21010
rect 29920 20946 29972 20952
rect 29932 20806 29960 20946
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 30378 6760 30434 6769
rect 30378 6695 30434 6704
rect 30392 6458 30420 6695
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30484 2650 30512 21490
rect 30932 10464 30984 10470
rect 30932 10406 30984 10412
rect 30944 9722 30972 10406
rect 30932 9716 30984 9722
rect 30932 9658 30984 9664
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 30760 3194 30788 8910
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30472 2644 30524 2650
rect 30472 2586 30524 2592
rect 31128 2514 31156 25434
rect 32324 21690 32352 37198
rect 33048 37120 33100 37126
rect 33048 37062 33100 37068
rect 33060 30326 33088 37062
rect 33140 36576 33192 36582
rect 33140 36518 33192 36524
rect 33048 30320 33100 30326
rect 33048 30262 33100 30268
rect 33152 30258 33180 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35452 34610 35480 37198
rect 35544 37126 35572 37318
rect 35992 37256 36044 37262
rect 35992 37198 36044 37204
rect 35532 37120 35584 37126
rect 35532 37062 35584 37068
rect 35532 36168 35584 36174
rect 35532 36110 35584 36116
rect 35440 34604 35492 34610
rect 35440 34546 35492 34552
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33232 32428 33284 32434
rect 33232 32370 33284 32376
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33244 29306 33272 32370
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 33692 30660 33744 30666
rect 33692 30602 33744 30608
rect 33232 29300 33284 29306
rect 33232 29242 33284 29248
rect 32404 26784 32456 26790
rect 32404 26726 32456 26732
rect 32312 21684 32364 21690
rect 32312 21626 32364 21632
rect 32416 21418 32444 26726
rect 32404 21412 32456 21418
rect 32404 21354 32456 21360
rect 31760 17196 31812 17202
rect 31760 17138 31812 17144
rect 31772 16590 31800 17138
rect 31760 16584 31812 16590
rect 31760 16526 31812 16532
rect 33048 10668 33100 10674
rect 33048 10610 33100 10616
rect 33060 8634 33088 10610
rect 33140 9988 33192 9994
rect 33140 9930 33192 9936
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 31390 8256 31446 8265
rect 31390 8191 31446 8200
rect 31404 8090 31432 8191
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31404 4622 31432 4762
rect 32312 4752 32364 4758
rect 32312 4694 32364 4700
rect 31392 4616 31444 4622
rect 31392 4558 31444 4564
rect 32324 2650 32352 4694
rect 33152 2650 33180 9930
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 33704 2446 33732 30602
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35452 28558 35480 34546
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34612 26512 34664 26518
rect 34612 26454 34664 26460
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34532 23322 34560 24754
rect 34624 23730 34652 26454
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34520 23316 34572 23322
rect 34520 23258 34572 23264
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35544 19922 35572 36110
rect 36004 35894 36032 37198
rect 36096 36854 36124 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 36084 36848 36136 36854
rect 36084 36790 36136 36796
rect 36176 36780 36228 36786
rect 36176 36722 36228 36728
rect 36188 36378 36216 36722
rect 37200 36378 37228 38791
rect 36176 36372 36228 36378
rect 36176 36314 36228 36320
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 36820 36168 36872 36174
rect 36820 36110 36872 36116
rect 37280 36168 37332 36174
rect 37280 36110 37332 36116
rect 35912 35866 36032 35894
rect 35912 29646 35940 35866
rect 36832 34746 36860 36110
rect 37292 35222 37320 36110
rect 37280 35216 37332 35222
rect 37280 35158 37332 35164
rect 37384 35086 37412 39200
rect 38106 37496 38162 37505
rect 38106 37431 38162 37440
rect 38120 36854 38148 37431
rect 38672 37330 38700 39200
rect 38660 37324 38712 37330
rect 38660 37266 38712 37272
rect 39316 36922 39344 39200
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 38108 36848 38160 36854
rect 38108 36790 38160 36796
rect 37924 36576 37976 36582
rect 37924 36518 37976 36524
rect 37832 35692 37884 35698
rect 37832 35634 37884 35640
rect 37372 35080 37424 35086
rect 37372 35022 37424 35028
rect 37464 34944 37516 34950
rect 37464 34886 37516 34892
rect 36820 34740 36872 34746
rect 36820 34682 36872 34688
rect 35992 34604 36044 34610
rect 35992 34546 36044 34552
rect 35900 29640 35952 29646
rect 35900 29582 35952 29588
rect 35900 27464 35952 27470
rect 35900 27406 35952 27412
rect 35912 25498 35940 27406
rect 36004 26586 36032 34546
rect 36452 32904 36504 32910
rect 36452 32846 36504 32852
rect 36464 28218 36492 32846
rect 37476 31346 37504 34886
rect 37464 31340 37516 31346
rect 37464 31282 37516 31288
rect 37004 30592 37056 30598
rect 37004 30534 37056 30540
rect 36452 28212 36504 28218
rect 36452 28154 36504 28160
rect 36084 27872 36136 27878
rect 36084 27814 36136 27820
rect 35992 26580 36044 26586
rect 35992 26522 36044 26528
rect 36096 26234 36124 27814
rect 37016 26994 37044 30534
rect 37740 29504 37792 29510
rect 37740 29446 37792 29452
rect 37004 26988 37056 26994
rect 37004 26930 37056 26936
rect 36004 26206 36124 26234
rect 35900 25492 35952 25498
rect 35900 25434 35952 25440
rect 36004 24750 36032 26206
rect 35992 24744 36044 24750
rect 35992 24686 36044 24692
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 36096 21146 36124 24142
rect 37752 23798 37780 29446
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37844 22794 37872 35634
rect 37752 22766 37872 22794
rect 36084 21140 36136 21146
rect 36084 21082 36136 21088
rect 37188 20936 37240 20942
rect 37188 20878 37240 20884
rect 37200 20505 37228 20878
rect 37752 20806 37780 22766
rect 37832 22636 37884 22642
rect 37832 22578 37884 22584
rect 37844 22234 37872 22578
rect 37832 22228 37884 22234
rect 37832 22170 37884 22176
rect 37832 20936 37884 20942
rect 37832 20878 37884 20884
rect 37740 20800 37792 20806
rect 37740 20742 37792 20748
rect 37186 20496 37242 20505
rect 37186 20431 37242 20440
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34440 18290 34468 19654
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34428 18284 34480 18290
rect 34428 18226 34480 18232
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35452 17338 35480 18226
rect 35440 17332 35492 17338
rect 35440 17274 35492 17280
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 36544 16108 36596 16114
rect 36544 16050 36596 16056
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 36556 14618 36584 16050
rect 37844 15026 37872 20878
rect 37936 16794 37964 36518
rect 38198 36136 38254 36145
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38200 32768 38252 32774
rect 38198 32736 38200 32745
rect 38252 32736 38254 32745
rect 38198 32671 38254 32680
rect 38200 32224 38252 32230
rect 38200 32166 38252 32172
rect 38212 32065 38240 32166
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38292 30728 38344 30734
rect 38290 30696 38292 30705
rect 38344 30696 38346 30705
rect 38290 30631 38346 30640
rect 38108 29572 38160 29578
rect 38108 29514 38160 29520
rect 38120 29345 38148 29514
rect 38106 29336 38162 29345
rect 38106 29271 38162 29280
rect 38292 28076 38344 28082
rect 38292 28018 38344 28024
rect 38304 27985 38332 28018
rect 38290 27976 38346 27985
rect 38290 27911 38346 27920
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38304 25945 38332 26318
rect 38290 25936 38346 25945
rect 38290 25871 38346 25880
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38200 24064 38252 24070
rect 38200 24006 38252 24012
rect 38212 23905 38240 24006
rect 38198 23896 38254 23905
rect 38198 23831 38254 23840
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38016 22432 38068 22438
rect 38016 22374 38068 22380
rect 38028 22030 38056 22374
rect 38016 22024 38068 22030
rect 38016 21966 38068 21972
rect 38016 21548 38068 21554
rect 38016 21490 38068 21496
rect 38028 18902 38056 21490
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 38304 19145 38332 19314
rect 38290 19136 38346 19145
rect 38290 19071 38346 19080
rect 38016 18896 38068 18902
rect 38016 18838 38068 18844
rect 38016 18080 38068 18086
rect 38016 18022 38068 18028
rect 38200 18080 38252 18086
rect 38200 18022 38252 18028
rect 37924 16788 37976 16794
rect 37924 16730 37976 16736
rect 38028 16590 38056 18022
rect 38212 17785 38240 18022
rect 38198 17776 38254 17785
rect 38198 17711 38254 17720
rect 38016 16584 38068 16590
rect 38016 16526 38068 16532
rect 38200 16448 38252 16454
rect 38198 16416 38200 16425
rect 38252 16416 38254 16425
rect 38198 16351 38254 16360
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 37832 15020 37884 15026
rect 37832 14962 37884 14968
rect 37924 14816 37976 14822
rect 37924 14758 37976 14764
rect 34520 14612 34572 14618
rect 34520 14554 34572 14560
rect 36544 14612 36596 14618
rect 36544 14554 36596 14560
rect 34532 10130 34560 14554
rect 34612 14408 34664 14414
rect 34612 14350 34664 14356
rect 37280 14408 37332 14414
rect 37280 14350 37332 14356
rect 34520 10124 34572 10130
rect 34520 10066 34572 10072
rect 34624 10010 34652 14350
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34808 13326 34836 14010
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 13320 34848 13326
rect 34796 13262 34848 13268
rect 37292 13258 37320 14350
rect 37280 13252 37332 13258
rect 37280 13194 37332 13200
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34440 9994 34652 10010
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 34428 9988 34652 9994
rect 34480 9982 34652 9988
rect 34428 9930 34480 9936
rect 37200 9625 37228 9998
rect 37186 9616 37242 9625
rect 37186 9551 37242 9560
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34428 8356 34480 8362
rect 34428 8298 34480 8304
rect 34440 7886 34468 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34060 6316 34112 6322
rect 34060 6258 34112 6264
rect 34072 4826 34100 6258
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34060 4820 34112 4826
rect 34060 4762 34112 4768
rect 34428 4480 34480 4486
rect 34428 4422 34480 4428
rect 34440 2446 34468 4422
rect 37188 4208 37240 4214
rect 37188 4150 37240 4156
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 34428 2440 34480 2446
rect 34428 2382 34480 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 28368 800 28396 2382
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29656 800 29684 2246
rect 30300 800 30328 2382
rect 31588 800 31616 2382
rect 32864 2372 32916 2378
rect 32864 2314 32916 2320
rect 32876 800 32904 2314
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 33520 800 33548 2246
rect 34808 800 34836 2246
rect 36096 800 36124 2246
rect 36740 800 36768 2382
rect 37200 1465 37228 4150
rect 37740 3732 37792 3738
rect 37740 3674 37792 3680
rect 37752 3058 37780 3674
rect 37936 3534 37964 14758
rect 38198 14376 38254 14385
rect 38198 14311 38254 14320
rect 38212 14278 38240 14311
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 38212 13025 38240 13126
rect 38198 13016 38254 13025
rect 38198 12951 38254 12960
rect 38292 12844 38344 12850
rect 38292 12786 38344 12792
rect 38108 12640 38160 12646
rect 38108 12582 38160 12588
rect 38120 12238 38148 12582
rect 38304 12345 38332 12786
rect 38290 12336 38346 12345
rect 38290 12271 38346 12280
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38108 11756 38160 11762
rect 38108 11698 38160 11704
rect 38120 11354 38148 11698
rect 38108 11348 38160 11354
rect 38108 11290 38160 11296
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38304 10985 38332 11086
rect 38290 10976 38346 10985
rect 38290 10911 38346 10920
rect 38108 10600 38160 10606
rect 38108 10542 38160 10548
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 38028 5234 38056 7686
rect 38120 6458 38148 10542
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38304 8265 38332 8434
rect 38290 8256 38346 8265
rect 38290 8191 38346 8200
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38346 7520
rect 38108 6452 38160 6458
rect 38108 6394 38160 6400
rect 38292 6316 38344 6322
rect 38292 6258 38344 6264
rect 38304 6225 38332 6258
rect 38290 6216 38346 6225
rect 38290 6151 38346 6160
rect 38016 5228 38068 5234
rect 38016 5170 38068 5176
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 38212 4865 38240 4966
rect 38198 4856 38254 4865
rect 38198 4791 38254 4800
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 38304 4185 38332 4558
rect 38290 4176 38346 4185
rect 38290 4111 38346 4120
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 32862 200 32918 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 36726 200 36782 800
rect 37476 785 37504 2926
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 37752 1834 37780 2382
rect 37740 1828 37792 1834
rect 37740 1770 37792 1776
rect 38028 800 38056 3334
rect 38212 2825 38240 3334
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 38198 2816 38254 2825
rect 38198 2751 38254 2760
rect 39316 800 39344 2926
rect 37462 776 37518 785
rect 37462 711 37518 720
rect 38014 200 38070 800
rect 39302 200 39358 800
rect 27988 128 28040 134
rect 27988 70 28040 76
rect 7196 60 7248 66
rect 7196 2 7248 8
rect 27344 60 27396 66
rect 27344 2 27396 8
<< via2 >>
rect 1582 38800 1638 38856
rect 1766 38120 1822 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2778 36760 2834 36816
rect 1582 35944 1638 36000
rect 1766 35436 1768 35456
rect 1768 35436 1820 35456
rect 1820 35436 1822 35456
rect 1766 35400 1822 35436
rect 1766 34720 1822 34776
rect 1766 33380 1822 33416
rect 1766 33360 1768 33380
rect 1768 33360 1820 33380
rect 1820 33360 1822 33380
rect 1582 32000 1638 32056
rect 1766 31320 1822 31376
rect 1766 29996 1768 30016
rect 1768 29996 1820 30016
rect 1820 29996 1822 30016
rect 1766 29960 1822 29996
rect 1766 28600 1822 28656
rect 1766 27276 1768 27296
rect 1768 27276 1820 27296
rect 1820 27276 1822 27296
rect 1766 27240 1822 27276
rect 1398 26560 1454 26616
rect 1122 12144 1178 12200
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1582 21800 1638 21856
rect 2318 26832 2374 26888
rect 1858 26560 1914 26616
rect 2134 23604 2136 23624
rect 2136 23604 2188 23624
rect 2188 23604 2190 23624
rect 2134 23568 2190 23604
rect 1858 17312 1914 17368
rect 1858 11872 1914 11928
rect 1766 8880 1822 8936
rect 1582 7520 1638 7576
rect 2502 24148 2504 24168
rect 2504 24148 2556 24168
rect 2556 24148 2558 24168
rect 2502 24112 2558 24148
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 2686 26324 2688 26344
rect 2688 26324 2740 26344
rect 2740 26324 2742 26344
rect 2686 26288 2742 26324
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 3238 26288 3294 26344
rect 2594 20576 2650 20632
rect 2226 13640 2282 13696
rect 2318 10804 2374 10840
rect 3974 25644 3976 25664
rect 3976 25644 4028 25664
rect 4028 25644 4030 25664
rect 3238 21936 3294 21992
rect 2962 20440 3018 20496
rect 2778 15680 2834 15736
rect 2870 11600 2926 11656
rect 2318 10784 2320 10804
rect 2320 10784 2372 10804
rect 2372 10784 2374 10804
rect 2778 10240 2834 10296
rect 2594 9172 2650 9208
rect 2594 9152 2596 9172
rect 2596 9152 2648 9172
rect 2648 9152 2650 9172
rect 1950 6316 2006 6352
rect 1950 6296 1952 6316
rect 1952 6296 2004 6316
rect 2004 6296 2006 6316
rect 1766 4120 1822 4176
rect 1582 3304 1638 3360
rect 3974 25608 4030 25644
rect 3974 24928 4030 24984
rect 3514 23196 3516 23216
rect 3516 23196 3568 23216
rect 3568 23196 3570 23216
rect 3514 23160 3570 23196
rect 3698 23024 3754 23080
rect 3330 18536 3386 18592
rect 3238 18400 3294 18456
rect 3330 17856 3386 17912
rect 3422 15272 3478 15328
rect 3330 14900 3332 14920
rect 3332 14900 3384 14920
rect 3384 14900 3386 14920
rect 3330 14864 3386 14900
rect 3330 12724 3332 12744
rect 3332 12724 3384 12744
rect 3384 12724 3386 12744
rect 3330 12688 3386 12724
rect 3882 22480 3938 22536
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 3882 21528 3938 21584
rect 3790 20712 3846 20768
rect 3606 19624 3662 19680
rect 3698 19508 3754 19544
rect 3698 19488 3700 19508
rect 3700 19488 3752 19508
rect 3752 19488 3754 19508
rect 3606 16904 3662 16960
rect 3790 17448 3846 17504
rect 3974 20576 4030 20632
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4434 21664 4490 21720
rect 4250 21392 4306 21448
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4986 24012 4988 24032
rect 4988 24012 5040 24032
rect 5040 24012 5042 24032
rect 4986 23976 5042 24012
rect 4894 23840 4950 23896
rect 4894 22480 4950 22536
rect 4526 20868 4582 20904
rect 4526 20848 4528 20868
rect 4528 20848 4580 20868
rect 4580 20848 4582 20868
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4342 19488 4398 19544
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3974 17720 4030 17776
rect 4526 17584 4582 17640
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 3790 16244 3846 16280
rect 3790 16224 3792 16244
rect 3792 16224 3844 16244
rect 3844 16224 3846 16244
rect 3238 12280 3294 12336
rect 3606 10512 3662 10568
rect 3238 9016 3294 9072
rect 2870 7928 2926 7984
rect 2686 5108 2688 5128
rect 2688 5108 2740 5128
rect 2740 5108 2742 5128
rect 2686 5072 2742 5108
rect 3606 6568 3662 6624
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12860 4068 12880
rect 4068 12860 4120 12880
rect 4120 12860 4122 12880
rect 4066 12824 4122 12860
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4250 12164 4306 12200
rect 4250 12144 4252 12164
rect 4252 12144 4304 12164
rect 4304 12144 4306 12164
rect 3974 12008 4030 12064
rect 5078 21800 5134 21856
rect 5354 23024 5410 23080
rect 5354 21664 5410 21720
rect 5170 18808 5226 18864
rect 4894 17076 4896 17096
rect 4896 17076 4948 17096
rect 4948 17076 4950 17096
rect 4894 17040 4950 17076
rect 4526 11736 4582 11792
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 9016 4122 9072
rect 3146 2624 3202 2680
rect 1766 2080 1822 2136
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4618 6160 4674 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4434 5244 4436 5264
rect 4436 5244 4488 5264
rect 4488 5244 4490 5264
rect 4434 5208 4490 5244
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4526 3984 4582 4040
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4342 3612 4344 3632
rect 4344 3612 4396 3632
rect 4396 3612 4398 3632
rect 4342 3576 4398 3612
rect 4066 3440 4122 3496
rect 4342 3476 4344 3496
rect 4344 3476 4396 3496
rect 4396 3476 4398 3496
rect 4342 3440 4398 3476
rect 3882 2488 3938 2544
rect 4802 7540 4858 7576
rect 4802 7520 4804 7540
rect 4804 7520 4856 7540
rect 4856 7520 4858 7540
rect 4710 4256 4766 4312
rect 5446 21256 5502 21312
rect 5446 17756 5448 17776
rect 5448 17756 5500 17776
rect 5500 17756 5502 17776
rect 5446 17720 5502 17756
rect 5446 17176 5502 17232
rect 5722 22480 5778 22536
rect 5722 21956 5778 21992
rect 5722 21936 5724 21956
rect 5724 21936 5776 21956
rect 5776 21936 5778 21956
rect 5722 21800 5778 21856
rect 5722 17992 5778 18048
rect 6458 26324 6460 26344
rect 6460 26324 6512 26344
rect 6512 26324 6514 26344
rect 6458 26288 6514 26324
rect 6090 23432 6146 23488
rect 5998 22752 6054 22808
rect 5906 22208 5962 22264
rect 5998 20304 6054 20360
rect 6182 22208 6238 22264
rect 6274 22072 6330 22128
rect 6274 21936 6330 21992
rect 6182 21004 6238 21040
rect 6182 20984 6184 21004
rect 6184 20984 6236 21004
rect 6236 20984 6238 21004
rect 6182 19780 6238 19816
rect 6182 19760 6184 19780
rect 6184 19760 6236 19780
rect 6236 19760 6238 19780
rect 6274 18536 6330 18592
rect 6090 17584 6146 17640
rect 5998 17312 6054 17368
rect 6550 21972 6552 21992
rect 6552 21972 6604 21992
rect 6604 21972 6606 21992
rect 6550 21936 6606 21972
rect 6458 20304 6514 20360
rect 7378 30368 7434 30424
rect 7010 23568 7066 23624
rect 6826 21392 6882 21448
rect 6734 20848 6790 20904
rect 6458 17312 6514 17368
rect 5538 13368 5594 13424
rect 5906 13368 5962 13424
rect 5722 13232 5778 13288
rect 5354 12180 5356 12200
rect 5356 12180 5408 12200
rect 5408 12180 5410 12200
rect 5354 12144 5410 12180
rect 5446 9696 5502 9752
rect 5906 11872 5962 11928
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3698 1536 3754 1592
rect 4066 2352 4122 2408
rect 5078 4276 5134 4312
rect 5078 4256 5080 4276
rect 5080 4256 5132 4276
rect 5132 4256 5134 4276
rect 5078 3984 5134 4040
rect 5078 3032 5134 3088
rect 5170 2896 5226 2952
rect 5722 5092 5778 5128
rect 5722 5072 5724 5092
rect 5724 5072 5776 5092
rect 5776 5072 5778 5092
rect 5722 4528 5778 4584
rect 6182 6840 6238 6896
rect 7010 20712 7066 20768
rect 7470 22072 7526 22128
rect 7010 19352 7066 19408
rect 6826 18808 6882 18864
rect 7102 19080 7158 19136
rect 7102 18536 7158 18592
rect 7010 18264 7066 18320
rect 6734 17040 6790 17096
rect 6826 12552 6882 12608
rect 8022 24112 8078 24168
rect 7470 19488 7526 19544
rect 7286 18944 7342 19000
rect 7194 16496 7250 16552
rect 7102 15020 7158 15056
rect 7102 15000 7104 15020
rect 7104 15000 7156 15020
rect 7156 15000 7158 15020
rect 7010 12416 7066 12472
rect 7654 16516 7710 16552
rect 7654 16496 7656 16516
rect 7656 16496 7708 16516
rect 7708 16496 7710 16516
rect 7654 16224 7710 16280
rect 7838 21800 7894 21856
rect 8114 18672 8170 18728
rect 8114 15544 8170 15600
rect 6826 10684 6828 10704
rect 6828 10684 6880 10704
rect 6880 10684 6882 10704
rect 6826 10648 6882 10684
rect 6550 9444 6606 9480
rect 6550 9424 6552 9444
rect 6552 9424 6604 9444
rect 6604 9424 6606 9444
rect 6734 8900 6790 8936
rect 6734 8880 6736 8900
rect 6736 8880 6788 8900
rect 6788 8880 6790 8900
rect 5814 3168 5870 3224
rect 6550 7248 6606 7304
rect 6918 5208 6974 5264
rect 6734 3984 6790 4040
rect 6550 3440 6606 3496
rect 6826 3576 6882 3632
rect 7470 12280 7526 12336
rect 7562 11348 7618 11384
rect 7562 11328 7564 11348
rect 7564 11328 7616 11348
rect 7616 11328 7618 11348
rect 7838 10104 7894 10160
rect 7194 6432 7250 6488
rect 7194 6024 7250 6080
rect 8298 22480 8354 22536
rect 8298 20868 8354 20904
rect 8298 20848 8300 20868
rect 8300 20848 8352 20868
rect 8352 20848 8354 20868
rect 8390 19488 8446 19544
rect 9770 30232 9826 30288
rect 9218 22480 9274 22536
rect 8390 15272 8446 15328
rect 8298 13232 8354 13288
rect 8850 18808 8906 18864
rect 8942 18536 8998 18592
rect 8758 15408 8814 15464
rect 8574 12416 8630 12472
rect 8482 10104 8538 10160
rect 7654 7112 7710 7168
rect 7378 4120 7434 4176
rect 7746 4936 7802 4992
rect 7838 3168 7894 3224
rect 8942 17740 8998 17776
rect 8942 17720 8944 17740
rect 8944 17720 8996 17740
rect 8996 17720 8998 17740
rect 8850 14456 8906 14512
rect 8850 13776 8906 13832
rect 8022 3168 8078 3224
rect 8574 8200 8630 8256
rect 9126 16632 9182 16688
rect 9954 21256 10010 21312
rect 9402 16904 9458 16960
rect 9862 19896 9918 19952
rect 9954 19388 9956 19408
rect 9956 19388 10008 19408
rect 10008 19388 10010 19408
rect 9954 19352 10010 19388
rect 9862 18400 9918 18456
rect 9770 17720 9826 17776
rect 9310 16788 9366 16824
rect 9310 16768 9312 16788
rect 9312 16768 9364 16788
rect 9364 16768 9366 16788
rect 9586 16768 9642 16824
rect 9310 16632 9366 16688
rect 9126 15272 9182 15328
rect 9586 16532 9588 16552
rect 9588 16532 9640 16552
rect 9640 16532 9642 16552
rect 9586 16496 9642 16532
rect 9310 15136 9366 15192
rect 9494 14340 9550 14376
rect 9494 14320 9496 14340
rect 9496 14320 9548 14340
rect 9548 14320 9550 14340
rect 9586 12960 9642 13016
rect 9310 11328 9366 11384
rect 8574 6840 8630 6896
rect 8574 6160 8630 6216
rect 7378 2896 7434 2952
rect 8850 7248 8906 7304
rect 8758 7112 8814 7168
rect 9770 16108 9826 16144
rect 9770 16088 9772 16108
rect 9772 16088 9824 16108
rect 9824 16088 9826 16108
rect 10230 18808 10286 18864
rect 10230 17448 10286 17504
rect 10782 22516 10784 22536
rect 10784 22516 10836 22536
rect 10836 22516 10838 22536
rect 10782 22480 10838 22516
rect 10506 21528 10562 21584
rect 10414 19216 10470 19272
rect 10506 16360 10562 16416
rect 10414 16224 10470 16280
rect 9678 11600 9734 11656
rect 10046 14048 10102 14104
rect 9954 11464 10010 11520
rect 10230 12960 10286 13016
rect 10230 12280 10286 12336
rect 10782 21956 10838 21992
rect 10782 21936 10784 21956
rect 10784 21936 10836 21956
rect 10836 21936 10838 21956
rect 10782 21664 10838 21720
rect 11058 21800 11114 21856
rect 10966 21004 11022 21040
rect 10966 20984 10968 21004
rect 10968 20984 11020 21004
rect 11020 20984 11022 21004
rect 11058 20712 11114 20768
rect 10966 19624 11022 19680
rect 10874 18808 10930 18864
rect 11058 18944 11114 19000
rect 10874 17856 10930 17912
rect 10874 17484 10876 17504
rect 10876 17484 10928 17504
rect 10928 17484 10930 17504
rect 10874 17448 10930 17484
rect 10874 16904 10930 16960
rect 10966 16632 11022 16688
rect 11518 21140 11574 21176
rect 11518 21120 11520 21140
rect 11520 21120 11572 21140
rect 11572 21120 11574 21140
rect 11426 20576 11482 20632
rect 11426 20032 11482 20088
rect 11518 19624 11574 19680
rect 10690 14356 10692 14376
rect 10692 14356 10744 14376
rect 10744 14356 10746 14376
rect 10690 14320 10746 14356
rect 10966 15816 11022 15872
rect 10598 12960 10654 13016
rect 10414 12280 10470 12336
rect 9678 9868 9680 9888
rect 9680 9868 9732 9888
rect 9732 9868 9734 9888
rect 9678 9832 9734 9868
rect 9218 8336 9274 8392
rect 9034 6840 9090 6896
rect 5262 1808 5318 1864
rect 6550 1944 6606 2000
rect 1398 720 1454 776
rect 9402 6740 9404 6760
rect 9404 6740 9456 6760
rect 9456 6740 9458 6760
rect 9402 6704 9458 6740
rect 9586 9596 9588 9616
rect 9588 9596 9640 9616
rect 9640 9596 9642 9616
rect 9586 9560 9642 9596
rect 10598 10920 10654 10976
rect 9678 8200 9734 8256
rect 9586 6976 9642 7032
rect 10414 8608 10470 8664
rect 9954 5480 10010 5536
rect 9862 5344 9918 5400
rect 9402 3884 9404 3904
rect 9404 3884 9456 3904
rect 9456 3884 9458 3904
rect 9402 3848 9458 3884
rect 10046 4664 10102 4720
rect 9678 2760 9734 2816
rect 10414 7792 10470 7848
rect 10874 9288 10930 9344
rect 10782 8880 10838 8936
rect 10230 3440 10286 3496
rect 10506 5752 10562 5808
rect 11426 18808 11482 18864
rect 11794 22208 11850 22264
rect 11794 21800 11850 21856
rect 11426 18536 11482 18592
rect 12070 18808 12126 18864
rect 12162 18708 12164 18728
rect 12164 18708 12216 18728
rect 12216 18708 12218 18728
rect 12162 18672 12218 18708
rect 11978 18572 11980 18592
rect 11980 18572 12032 18592
rect 12032 18572 12034 18592
rect 11978 18536 12034 18572
rect 11886 17720 11942 17776
rect 11334 15680 11390 15736
rect 11150 14592 11206 14648
rect 11150 12588 11152 12608
rect 11152 12588 11204 12608
rect 11204 12588 11206 12608
rect 11150 12552 11206 12588
rect 11150 11872 11206 11928
rect 11242 11056 11298 11112
rect 11610 16632 11666 16688
rect 12070 17992 12126 18048
rect 12438 19216 12494 19272
rect 12714 19660 12716 19680
rect 12716 19660 12768 19680
rect 12768 19660 12770 19680
rect 12714 19624 12770 19660
rect 12346 18400 12402 18456
rect 11702 16088 11758 16144
rect 11426 13232 11482 13288
rect 11702 14184 11758 14240
rect 12346 16768 12402 16824
rect 12070 16088 12126 16144
rect 12070 14592 12126 14648
rect 11518 12688 11574 12744
rect 11794 12008 11850 12064
rect 10966 8064 11022 8120
rect 11334 10784 11390 10840
rect 11150 7656 11206 7712
rect 11150 7520 11206 7576
rect 10966 7384 11022 7440
rect 11058 7248 11114 7304
rect 10874 5616 10930 5672
rect 10598 2760 10654 2816
rect 12346 15544 12402 15600
rect 12990 18264 13046 18320
rect 12254 15136 12310 15192
rect 12530 15136 12586 15192
rect 12070 12280 12126 12336
rect 13358 23432 13414 23488
rect 13358 22208 13414 22264
rect 13266 21972 13268 21992
rect 13268 21972 13320 21992
rect 13320 21972 13322 21992
rect 13266 21936 13322 21972
rect 13358 20304 13414 20360
rect 14830 23724 14886 23760
rect 14830 23704 14832 23724
rect 14832 23704 14884 23724
rect 14884 23704 14886 23724
rect 14186 21548 14242 21584
rect 14186 21528 14188 21548
rect 14188 21528 14240 21548
rect 14240 21528 14242 21548
rect 13450 18536 13506 18592
rect 13450 18128 13506 18184
rect 13358 16224 13414 16280
rect 13174 12688 13230 12744
rect 11610 9968 11666 10024
rect 11518 9424 11574 9480
rect 11886 10140 11888 10160
rect 11888 10140 11940 10160
rect 11940 10140 11942 10160
rect 11886 10104 11942 10140
rect 12162 9988 12218 10024
rect 12162 9968 12164 9988
rect 12164 9968 12216 9988
rect 12216 9968 12218 9988
rect 11518 8880 11574 8936
rect 11794 9152 11850 9208
rect 12530 9152 12586 9208
rect 12162 8200 12218 8256
rect 12070 7656 12126 7712
rect 11150 4256 11206 4312
rect 12070 5208 12126 5264
rect 11518 3848 11574 3904
rect 11978 5072 12034 5128
rect 12254 5480 12310 5536
rect 12346 5208 12402 5264
rect 12162 4528 12218 4584
rect 12070 4392 12126 4448
rect 12162 3848 12218 3904
rect 11978 3476 11980 3496
rect 11980 3476 12032 3496
rect 12032 3476 12034 3496
rect 11978 3440 12034 3476
rect 12622 6024 12678 6080
rect 12622 5616 12678 5672
rect 12346 4392 12402 4448
rect 12530 4528 12586 4584
rect 13082 10920 13138 10976
rect 12898 6432 12954 6488
rect 13358 15852 13360 15872
rect 13360 15852 13412 15872
rect 13412 15852 13414 15872
rect 13358 15816 13414 15852
rect 13358 15544 13414 15600
rect 13634 17312 13690 17368
rect 14002 19352 14058 19408
rect 13818 18400 13874 18456
rect 13818 17484 13820 17504
rect 13820 17484 13872 17504
rect 13872 17484 13874 17504
rect 13818 17448 13874 17484
rect 13726 17176 13782 17232
rect 13818 16632 13874 16688
rect 13450 12552 13506 12608
rect 13266 8744 13322 8800
rect 13634 11872 13690 11928
rect 14370 20304 14426 20360
rect 14186 18536 14242 18592
rect 14094 16360 14150 16416
rect 14278 15816 14334 15872
rect 14278 13640 14334 13696
rect 13818 10784 13874 10840
rect 13266 5888 13322 5944
rect 13266 5616 13322 5672
rect 13542 6160 13598 6216
rect 13542 5752 13598 5808
rect 13542 4392 13598 4448
rect 13450 3984 13506 4040
rect 14094 12008 14150 12064
rect 14462 19624 14518 19680
rect 14554 18264 14610 18320
rect 14278 12688 14334 12744
rect 14278 10104 14334 10160
rect 14186 8744 14242 8800
rect 14094 8608 14150 8664
rect 14002 7792 14058 7848
rect 13910 5480 13966 5536
rect 14278 6568 14334 6624
rect 14094 4936 14150 4992
rect 14002 4800 14058 4856
rect 14278 4548 14334 4584
rect 14278 4528 14280 4548
rect 14280 4528 14332 4548
rect 14332 4528 14334 4548
rect 13910 3984 13966 4040
rect 14186 3712 14242 3768
rect 14094 1672 14150 1728
rect 14922 21936 14978 21992
rect 15014 20440 15070 20496
rect 15014 18148 15070 18184
rect 15014 18128 15016 18148
rect 15016 18128 15068 18148
rect 15068 18128 15070 18148
rect 15014 15036 15016 15056
rect 15016 15036 15068 15056
rect 15068 15036 15070 15056
rect 15014 15000 15070 15036
rect 15290 20712 15346 20768
rect 15474 19760 15530 19816
rect 15382 19488 15438 19544
rect 15290 17720 15346 17776
rect 15382 17448 15438 17504
rect 15290 16224 15346 16280
rect 15934 22208 15990 22264
rect 16026 22072 16082 22128
rect 15842 20440 15898 20496
rect 15658 20340 15660 20360
rect 15660 20340 15712 20360
rect 15712 20340 15714 20360
rect 15658 20304 15714 20340
rect 15658 19896 15714 19952
rect 15566 15680 15622 15736
rect 15474 15136 15530 15192
rect 14922 12960 14978 13016
rect 14554 8064 14610 8120
rect 14646 6840 14702 6896
rect 14370 3576 14426 3632
rect 14462 2896 14518 2952
rect 15106 12552 15162 12608
rect 15014 8880 15070 8936
rect 15198 12008 15254 12064
rect 14922 6432 14978 6488
rect 15014 3848 15070 3904
rect 15474 11328 15530 11384
rect 16578 20984 16634 21040
rect 15750 13368 15806 13424
rect 15658 12724 15660 12744
rect 15660 12724 15712 12744
rect 15712 12724 15714 12744
rect 15658 12688 15714 12724
rect 15474 7520 15530 7576
rect 15290 5616 15346 5672
rect 15382 5344 15438 5400
rect 15198 3304 15254 3360
rect 15382 4120 15438 4176
rect 15750 9152 15806 9208
rect 16118 16788 16174 16824
rect 16118 16768 16120 16788
rect 16120 16768 16172 16788
rect 16172 16768 16174 16788
rect 16118 14864 16174 14920
rect 16118 12960 16174 13016
rect 16026 12316 16028 12336
rect 16028 12316 16080 12336
rect 16080 12316 16082 12336
rect 16026 12280 16082 12316
rect 16578 16904 16634 16960
rect 17314 22888 17370 22944
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 17774 23432 17830 23488
rect 17498 21256 17554 21312
rect 17130 20032 17186 20088
rect 16854 17992 16910 18048
rect 15934 9424 15990 9480
rect 17130 15308 17132 15328
rect 17132 15308 17184 15328
rect 17184 15308 17186 15328
rect 17130 15272 17186 15308
rect 17038 13232 17094 13288
rect 17038 12688 17094 12744
rect 16670 11464 16726 11520
rect 16578 10104 16634 10160
rect 16118 6704 16174 6760
rect 16118 6160 16174 6216
rect 16026 5516 16028 5536
rect 16028 5516 16080 5536
rect 16080 5516 16082 5536
rect 16026 5480 16082 5516
rect 15750 4120 15806 4176
rect 15842 3576 15898 3632
rect 16026 4392 16082 4448
rect 14922 2760 14978 2816
rect 15382 2624 15438 2680
rect 16026 3188 16082 3224
rect 16026 3168 16028 3188
rect 16028 3168 16080 3188
rect 16080 3168 16082 3188
rect 16578 8064 16634 8120
rect 16578 6976 16634 7032
rect 16302 6704 16358 6760
rect 16486 5888 16542 5944
rect 16578 5752 16634 5808
rect 16486 3576 16542 3632
rect 16394 3304 16450 3360
rect 17222 11192 17278 11248
rect 17038 10648 17094 10704
rect 16762 6840 16818 6896
rect 17682 21664 17738 21720
rect 17866 17856 17922 17912
rect 17590 15000 17646 15056
rect 18326 21800 18382 21856
rect 18602 19796 18604 19816
rect 18604 19796 18656 19816
rect 18656 19796 18658 19816
rect 18602 19760 18658 19796
rect 17314 8608 17370 8664
rect 17130 8200 17186 8256
rect 17590 8336 17646 8392
rect 18142 14048 18198 14104
rect 17958 13504 18014 13560
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19430 23432 19486 23488
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19246 18400 19302 18456
rect 18142 12280 18198 12336
rect 18050 11328 18106 11384
rect 17774 8916 17776 8936
rect 17776 8916 17828 8936
rect 17828 8916 17830 8936
rect 17774 8880 17830 8916
rect 18142 8744 18198 8800
rect 17406 5344 17462 5400
rect 17406 4936 17462 4992
rect 17314 4800 17370 4856
rect 17222 2624 17278 2680
rect 17682 7520 17738 7576
rect 17590 6568 17646 6624
rect 17590 5208 17646 5264
rect 17958 7692 17960 7712
rect 17960 7692 18012 7712
rect 18012 7692 18014 7712
rect 17958 7656 18014 7692
rect 17774 4936 17830 4992
rect 17682 4820 17738 4856
rect 17682 4800 17684 4820
rect 17684 4800 17736 4820
rect 17736 4800 17738 4820
rect 17682 4120 17738 4176
rect 17682 3848 17738 3904
rect 18694 10920 18750 10976
rect 18970 9832 19026 9888
rect 18694 8608 18750 8664
rect 18326 4256 18382 4312
rect 18694 6704 18750 6760
rect 18510 6568 18566 6624
rect 18878 8780 18880 8800
rect 18880 8780 18932 8800
rect 18932 8780 18934 8800
rect 18878 8744 18934 8780
rect 19062 8608 19118 8664
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19798 21428 19800 21448
rect 19800 21428 19852 21448
rect 19852 21428 19854 21448
rect 19798 21392 19854 21428
rect 20166 20848 20222 20904
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 20166 17176 20222 17232
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19614 12724 19616 12744
rect 19616 12724 19668 12744
rect 19668 12724 19670 12744
rect 19614 12688 19670 12724
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19982 11056 20038 11112
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19982 10784 20038 10840
rect 19338 10648 19394 10704
rect 19706 10376 19762 10432
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19982 9696 20038 9752
rect 19338 8880 19394 8936
rect 19338 8780 19340 8800
rect 19340 8780 19392 8800
rect 19392 8780 19394 8800
rect 19338 8744 19394 8780
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19982 8608 20038 8664
rect 20258 10376 20314 10432
rect 20166 8744 20222 8800
rect 20258 8336 20314 8392
rect 19890 7792 19946 7848
rect 20074 7828 20076 7848
rect 20076 7828 20128 7848
rect 20128 7828 20130 7848
rect 20074 7792 20130 7828
rect 19982 7656 20038 7712
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 18694 5652 18696 5672
rect 18696 5652 18748 5672
rect 18748 5652 18750 5672
rect 18694 5616 18750 5652
rect 19338 6740 19340 6760
rect 19340 6740 19392 6760
rect 19392 6740 19394 6760
rect 19338 6704 19394 6740
rect 19154 5480 19210 5536
rect 19246 5344 19302 5400
rect 19154 4936 19210 4992
rect 19982 6568 20038 6624
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19522 5652 19524 5672
rect 19524 5652 19576 5672
rect 19576 5652 19578 5672
rect 19522 5616 19578 5652
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 20442 7656 20498 7712
rect 21086 12552 21142 12608
rect 21270 15408 21326 15464
rect 20994 10412 20996 10432
rect 20996 10412 21048 10432
rect 21048 10412 21050 10432
rect 20994 10376 21050 10412
rect 21270 9968 21326 10024
rect 20350 7384 20406 7440
rect 20166 5344 20222 5400
rect 19430 4936 19486 4992
rect 20442 5480 20498 5536
rect 20902 5344 20958 5400
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19338 4120 19394 4176
rect 20166 4256 20222 4312
rect 20442 4528 20498 4584
rect 20534 3984 20590 4040
rect 20718 4120 20774 4176
rect 19062 2760 19118 2816
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20074 3340 20076 3360
rect 20076 3340 20128 3360
rect 20128 3340 20130 3360
rect 20074 3304 20130 3340
rect 20166 3168 20222 3224
rect 19614 3052 19670 3088
rect 19614 3032 19616 3052
rect 19616 3032 19668 3052
rect 19668 3032 19670 3052
rect 19982 3032 20038 3088
rect 20902 4256 20958 4312
rect 20534 3304 20590 3360
rect 20718 3304 20774 3360
rect 20166 2896 20222 2952
rect 20350 2896 20406 2952
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21914 11076 21970 11112
rect 21914 11056 21916 11076
rect 21916 11056 21968 11076
rect 21968 11056 21970 11076
rect 21546 10668 21602 10704
rect 21546 10648 21548 10668
rect 21548 10648 21600 10668
rect 21600 10648 21602 10668
rect 22098 10376 22154 10432
rect 21822 9988 21878 10024
rect 21822 9968 21824 9988
rect 21824 9968 21876 9988
rect 21876 9968 21878 9988
rect 22558 11600 22614 11656
rect 23846 17040 23902 17096
rect 23202 14456 23258 14512
rect 21270 5888 21326 5944
rect 21178 5752 21234 5808
rect 21362 5752 21418 5808
rect 21730 8336 21786 8392
rect 22006 8492 22062 8528
rect 22006 8472 22008 8492
rect 22008 8472 22060 8492
rect 22060 8472 22062 8492
rect 22834 9696 22890 9752
rect 22466 8064 22522 8120
rect 22374 7792 22430 7848
rect 22006 6976 22062 7032
rect 21822 6024 21878 6080
rect 21270 5344 21326 5400
rect 21086 5072 21142 5128
rect 21638 5616 21694 5672
rect 21822 5616 21878 5672
rect 21730 5344 21786 5400
rect 21822 3576 21878 3632
rect 22098 5480 22154 5536
rect 22006 4936 22062 4992
rect 22006 4700 22008 4720
rect 22008 4700 22060 4720
rect 22060 4700 22062 4720
rect 22006 4664 22062 4700
rect 22098 3612 22100 3632
rect 22100 3612 22152 3632
rect 22152 3612 22154 3632
rect 22098 3576 22154 3612
rect 21914 2896 21970 2952
rect 21638 2760 21694 2816
rect 22098 1808 22154 1864
rect 22466 3032 22522 3088
rect 23570 13232 23626 13288
rect 23386 12860 23388 12880
rect 23388 12860 23440 12880
rect 23440 12860 23442 12880
rect 23386 12824 23442 12860
rect 23294 12436 23350 12472
rect 23294 12416 23296 12436
rect 23296 12416 23348 12436
rect 23348 12416 23350 12436
rect 23294 11736 23350 11792
rect 23294 10512 23350 10568
rect 23110 9152 23166 9208
rect 22926 7384 22982 7440
rect 22742 5072 22798 5128
rect 22742 4276 22798 4312
rect 22742 4256 22744 4276
rect 22744 4256 22796 4276
rect 22796 4256 22798 4276
rect 22834 3848 22890 3904
rect 22650 3168 22706 3224
rect 22558 2760 22614 2816
rect 23662 10240 23718 10296
rect 23386 9288 23442 9344
rect 23570 6160 23626 6216
rect 23294 5616 23350 5672
rect 23386 4800 23442 4856
rect 23662 4548 23718 4584
rect 23662 4528 23664 4548
rect 23664 4528 23716 4548
rect 23716 4528 23718 4548
rect 23846 9988 23902 10024
rect 23846 9968 23848 9988
rect 23848 9968 23900 9988
rect 23900 9968 23902 9988
rect 24122 10804 24178 10840
rect 24122 10784 24124 10804
rect 24124 10784 24176 10804
rect 24176 10784 24178 10804
rect 23846 9424 23902 9480
rect 23846 7520 23902 7576
rect 23938 6568 23994 6624
rect 23294 3712 23350 3768
rect 22742 2624 22798 2680
rect 23386 2488 23442 2544
rect 23386 2352 23442 2408
rect 23938 1672 23994 1728
rect 24398 21392 24454 21448
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 25134 19080 25190 19136
rect 25686 19080 25742 19136
rect 24674 14592 24730 14648
rect 24398 9560 24454 9616
rect 24858 12144 24914 12200
rect 25042 10104 25098 10160
rect 27618 16108 27674 16144
rect 27618 16088 27620 16108
rect 27620 16088 27672 16108
rect 27672 16088 27674 16108
rect 25226 9016 25282 9072
rect 25318 8608 25374 8664
rect 24674 6296 24730 6352
rect 25226 7928 25282 7984
rect 24858 7284 24860 7304
rect 24860 7284 24912 7304
rect 24912 7284 24914 7304
rect 24858 7248 24914 7284
rect 24858 7112 24914 7168
rect 24030 1536 24086 1592
rect 25502 4392 25558 4448
rect 25870 5208 25926 5264
rect 26054 6840 26110 6896
rect 27342 11056 27398 11112
rect 28170 5752 28226 5808
rect 26606 3340 26608 3360
rect 26608 3340 26660 3360
rect 26660 3340 26662 3360
rect 26606 3304 26662 3340
rect 27158 1944 27214 2000
rect 27986 3576 28042 3632
rect 27802 3440 27858 3496
rect 30378 6704 30434 6760
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 31390 8200 31446 8256
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 37186 38800 37242 38856
rect 38106 37440 38162 37496
rect 37186 20440 37242 20496
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38198 36080 38254 36136
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 34040 38254 34096
rect 38198 32716 38200 32736
rect 38200 32716 38252 32736
rect 38252 32716 38254 32736
rect 38198 32680 38254 32716
rect 38198 32000 38254 32056
rect 38290 30676 38292 30696
rect 38292 30676 38344 30696
rect 38344 30676 38346 30696
rect 38290 30640 38346 30676
rect 38106 29280 38162 29336
rect 38290 27920 38346 27976
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38290 25880 38346 25936
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38198 23840 38254 23896
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 21120 38254 21176
rect 38290 19080 38346 19136
rect 38198 17720 38254 17776
rect 38198 16396 38200 16416
rect 38200 16396 38252 16416
rect 38252 16396 38254 16416
rect 38198 16360 38254 16396
rect 38198 15680 38254 15736
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 37186 9560 37242 9616
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38198 14320 38254 14376
rect 38198 12960 38254 13016
rect 38290 12280 38346 12336
rect 38290 10920 38346 10976
rect 38290 8200 38346 8256
rect 38290 7520 38346 7576
rect 38290 6160 38346 6216
rect 38198 4800 38254 4856
rect 38290 4120 38346 4176
rect 37186 1400 37242 1456
rect 38198 2760 38254 2816
rect 37462 720 37518 776
<< metal3 >>
rect 200 38858 800 38888
rect 1577 38858 1643 38861
rect 200 38856 1643 38858
rect 200 38800 1582 38856
rect 1638 38800 1643 38856
rect 200 38798 1643 38800
rect 200 38768 800 38798
rect 1577 38795 1643 38798
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 200 38178 800 38208
rect 1761 38178 1827 38181
rect 200 38176 1827 38178
rect 200 38120 1766 38176
rect 1822 38120 1827 38176
rect 200 38118 1827 38120
rect 200 38088 800 38118
rect 1761 38115 1827 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 38101 37498 38167 37501
rect 39200 37498 39800 37528
rect 38101 37496 39800 37498
rect 38101 37440 38106 37496
rect 38162 37440 39800 37496
rect 38101 37438 39800 37440
rect 38101 37435 38167 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 2773 36818 2839 36821
rect 200 36816 2839 36818
rect 200 36760 2778 36816
rect 2834 36760 2839 36816
rect 200 36758 2839 36760
rect 200 36728 800 36758
rect 2773 36755 2839 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 1577 36002 1643 36005
rect 2446 36002 2452 36004
rect 1577 36000 2452 36002
rect 1577 35944 1582 36000
rect 1638 35944 2452 36000
rect 1577 35942 2452 35944
rect 1577 35939 1643 35942
rect 2446 35940 2452 35942
rect 2516 35940 2522 36004
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35458 800 35488
rect 1761 35458 1827 35461
rect 200 35456 1827 35458
rect 200 35400 1766 35456
rect 1822 35400 1827 35456
rect 200 35398 1827 35400
rect 200 35368 800 35398
rect 1761 35395 1827 35398
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 200 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1761 34778 1827 34781
rect 200 34776 1827 34778
rect 200 34720 1766 34776
rect 1822 34720 1827 34776
rect 200 34718 1827 34720
rect 200 34688 800 34718
rect 1761 34715 1827 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 38193 32738 38259 32741
rect 39200 32738 39800 32768
rect 38193 32736 39800 32738
rect 38193 32680 38198 32736
rect 38254 32680 39800 32736
rect 38193 32678 39800 32680
rect 38193 32675 38259 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31968 800 31998
rect 1577 31995 1643 31998
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 200 31378 800 31408
rect 1761 31378 1827 31381
rect 200 31376 1827 31378
rect 200 31320 1766 31376
rect 1822 31320 1827 31376
rect 200 31318 1827 31320
rect 200 31288 800 31318
rect 1761 31315 1827 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 38285 30698 38351 30701
rect 39200 30698 39800 30728
rect 38285 30696 39800 30698
rect 38285 30640 38290 30696
rect 38346 30640 39800 30696
rect 38285 30638 39800 30640
rect 38285 30635 38351 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 6126 30364 6132 30428
rect 6196 30426 6202 30428
rect 7373 30426 7439 30429
rect 6196 30424 7439 30426
rect 6196 30368 7378 30424
rect 7434 30368 7439 30424
rect 6196 30366 7439 30368
rect 6196 30364 6202 30366
rect 7373 30363 7439 30366
rect 9765 30290 9831 30293
rect 18086 30290 18092 30292
rect 9765 30288 18092 30290
rect 9765 30232 9770 30288
rect 9826 30232 18092 30288
rect 9765 30230 18092 30232
rect 9765 30227 9831 30230
rect 18086 30228 18092 30230
rect 18156 30228 18162 30292
rect 200 30018 800 30048
rect 1761 30018 1827 30021
rect 200 30016 1827 30018
rect 200 29960 1766 30016
rect 1822 29960 1827 30016
rect 200 29958 1827 29960
rect 200 29928 800 29958
rect 1761 29955 1827 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 38101 29338 38167 29341
rect 39200 29338 39800 29368
rect 38101 29336 39800 29338
rect 38101 29280 38106 29336
rect 38162 29280 39800 29336
rect 38101 29278 39800 29280
rect 38101 29275 38167 29278
rect 39200 29248 39800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 38285 27978 38351 27981
rect 39200 27978 39800 28008
rect 38285 27976 39800 27978
rect 38285 27920 38290 27976
rect 38346 27920 39800 27976
rect 38285 27918 39800 27920
rect 38285 27915 38351 27918
rect 39200 27888 39800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 1710 26828 1716 26892
rect 1780 26890 1786 26892
rect 2313 26890 2379 26893
rect 1780 26888 2379 26890
rect 1780 26832 2318 26888
rect 2374 26832 2379 26888
rect 1780 26830 2379 26832
rect 1780 26828 1786 26830
rect 2313 26827 2379 26830
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1393 26618 1459 26621
rect 200 26616 1459 26618
rect 200 26560 1398 26616
rect 1454 26560 1459 26616
rect 200 26558 1459 26560
rect 200 26528 800 26558
rect 1393 26555 1459 26558
rect 1853 26618 1919 26621
rect 2630 26618 2636 26620
rect 1853 26616 2636 26618
rect 1853 26560 1858 26616
rect 1914 26560 2636 26616
rect 1853 26558 2636 26560
rect 1853 26555 1919 26558
rect 2630 26556 2636 26558
rect 2700 26556 2706 26620
rect 1894 26284 1900 26348
rect 1964 26346 1970 26348
rect 2681 26346 2747 26349
rect 1964 26344 2747 26346
rect 1964 26288 2686 26344
rect 2742 26288 2747 26344
rect 1964 26286 2747 26288
rect 1964 26284 1970 26286
rect 2681 26283 2747 26286
rect 3233 26346 3299 26349
rect 6453 26348 6519 26349
rect 3366 26346 3372 26348
rect 3233 26344 3372 26346
rect 3233 26288 3238 26344
rect 3294 26288 3372 26344
rect 3233 26286 3372 26288
rect 3233 26283 3299 26286
rect 3366 26284 3372 26286
rect 3436 26284 3442 26348
rect 6453 26346 6500 26348
rect 6408 26344 6500 26346
rect 6408 26288 6458 26344
rect 6408 26286 6500 26288
rect 6453 26284 6500 26286
rect 6564 26284 6570 26348
rect 6453 26283 6519 26284
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 3734 25604 3740 25668
rect 3804 25666 3810 25668
rect 3969 25666 4035 25669
rect 3804 25664 4035 25666
rect 3804 25608 3974 25664
rect 4030 25608 4035 25664
rect 3804 25606 4035 25608
rect 3804 25604 3810 25606
rect 3969 25603 4035 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25168 800 25198
rect 1577 25195 1643 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 3969 24988 4035 24989
rect 3918 24986 3924 24988
rect 3878 24926 3924 24986
rect 3988 24984 4035 24988
rect 4030 24928 4035 24984
rect 3918 24924 3924 24926
rect 3988 24924 4035 24928
rect 3969 24923 4035 24924
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 2497 24170 2563 24173
rect 8017 24170 8083 24173
rect 2497 24168 8083 24170
rect 2497 24112 2502 24168
rect 2558 24112 8022 24168
rect 8078 24112 8083 24168
rect 2497 24110 8083 24112
rect 2497 24107 2563 24110
rect 8017 24107 8083 24110
rect 4654 23972 4660 24036
rect 4724 24034 4730 24036
rect 4981 24034 5047 24037
rect 4724 24032 5047 24034
rect 4724 23976 4986 24032
rect 5042 23976 5047 24032
rect 4724 23974 5047 23976
rect 4724 23972 4730 23974
rect 4981 23971 5047 23974
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4889 23898 4955 23901
rect 10726 23898 10732 23900
rect 200 23896 4955 23898
rect 200 23840 4894 23896
rect 4950 23840 4955 23896
rect 200 23838 4955 23840
rect 200 23808 800 23838
rect 4889 23835 4955 23838
rect 5398 23838 10732 23898
rect 2129 23626 2195 23629
rect 5398 23626 5458 23838
rect 10726 23836 10732 23838
rect 10796 23836 10802 23900
rect 38193 23898 38259 23901
rect 39200 23898 39800 23928
rect 38193 23896 39800 23898
rect 38193 23840 38198 23896
rect 38254 23840 39800 23896
rect 38193 23838 39800 23840
rect 38193 23835 38259 23838
rect 39200 23808 39800 23838
rect 5574 23700 5580 23764
rect 5644 23762 5650 23764
rect 14825 23762 14891 23765
rect 5644 23760 14891 23762
rect 5644 23704 14830 23760
rect 14886 23704 14891 23760
rect 5644 23702 14891 23704
rect 5644 23700 5650 23702
rect 14825 23699 14891 23702
rect 2129 23624 5458 23626
rect 2129 23568 2134 23624
rect 2190 23568 5458 23624
rect 2129 23566 5458 23568
rect 7005 23626 7071 23629
rect 7230 23626 7236 23628
rect 7005 23624 7236 23626
rect 7005 23568 7010 23624
rect 7066 23568 7236 23624
rect 7005 23566 7236 23568
rect 2129 23563 2195 23566
rect 7005 23563 7071 23566
rect 7230 23564 7236 23566
rect 7300 23564 7306 23628
rect 6085 23490 6151 23493
rect 11094 23490 11100 23492
rect 6085 23488 11100 23490
rect 6085 23432 6090 23488
rect 6146 23432 11100 23488
rect 6085 23430 11100 23432
rect 6085 23427 6151 23430
rect 11094 23428 11100 23430
rect 11164 23428 11170 23492
rect 12566 23428 12572 23492
rect 12636 23490 12642 23492
rect 13353 23490 13419 23493
rect 12636 23488 13419 23490
rect 12636 23432 13358 23488
rect 13414 23432 13419 23488
rect 12636 23430 13419 23432
rect 12636 23428 12642 23430
rect 13353 23427 13419 23430
rect 17769 23490 17835 23493
rect 19425 23490 19491 23493
rect 17769 23488 19491 23490
rect 17769 23432 17774 23488
rect 17830 23432 19430 23488
rect 19486 23432 19491 23488
rect 17769 23430 19491 23432
rect 17769 23427 17835 23430
rect 19425 23427 19491 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 3509 23218 3575 23221
rect 200 23216 3575 23218
rect 200 23160 3514 23216
rect 3570 23160 3575 23216
rect 200 23158 3575 23160
rect 200 23128 800 23158
rect 3509 23155 3575 23158
rect 3693 23082 3759 23085
rect 5349 23082 5415 23085
rect 3693 23080 5415 23082
rect 3693 23024 3698 23080
rect 3754 23024 5354 23080
rect 5410 23024 5415 23080
rect 3693 23022 5415 23024
rect 3693 23019 3759 23022
rect 5349 23019 5415 23022
rect 15510 22884 15516 22948
rect 15580 22946 15586 22948
rect 17309 22946 17375 22949
rect 15580 22944 17375 22946
rect 15580 22888 17314 22944
rect 17370 22888 17375 22944
rect 15580 22886 17375 22888
rect 15580 22884 15586 22886
rect 17309 22883 17375 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 5993 22812 6059 22813
rect 5942 22810 5948 22812
rect 5902 22750 5948 22810
rect 6012 22808 6059 22812
rect 6054 22752 6059 22808
rect 5942 22748 5948 22750
rect 6012 22748 6059 22752
rect 5993 22747 6059 22748
rect 2814 22612 2820 22676
rect 2884 22674 2890 22676
rect 15510 22674 15516 22676
rect 2884 22614 15516 22674
rect 2884 22612 2890 22614
rect 15510 22612 15516 22614
rect 15580 22612 15586 22676
rect 3877 22538 3943 22541
rect 4889 22538 4955 22541
rect 5717 22540 5783 22541
rect 5717 22538 5764 22540
rect 3877 22536 4955 22538
rect 3877 22480 3882 22536
rect 3938 22480 4894 22536
rect 4950 22480 4955 22536
rect 3877 22478 4955 22480
rect 5672 22536 5764 22538
rect 5828 22538 5834 22540
rect 8293 22538 8359 22541
rect 5828 22536 8359 22538
rect 5672 22480 5722 22536
rect 5828 22480 8298 22536
rect 8354 22480 8359 22536
rect 5672 22478 5764 22480
rect 3877 22475 3943 22478
rect 4889 22475 4955 22478
rect 5717 22476 5764 22478
rect 5828 22478 8359 22480
rect 5828 22476 5834 22478
rect 5717 22475 5783 22476
rect 8293 22475 8359 22478
rect 9213 22538 9279 22541
rect 10777 22538 10843 22541
rect 9213 22536 10843 22538
rect 9213 22480 9218 22536
rect 9274 22480 10782 22536
rect 10838 22480 10843 22536
rect 9213 22478 10843 22480
rect 9213 22475 9279 22478
rect 10777 22475 10843 22478
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 5901 22266 5967 22269
rect 6177 22266 6243 22269
rect 5901 22264 6243 22266
rect 5901 22208 5906 22264
rect 5962 22208 6182 22264
rect 6238 22208 6243 22264
rect 5901 22206 6243 22208
rect 5901 22203 5967 22206
rect 6177 22203 6243 22206
rect 11789 22266 11855 22269
rect 13353 22266 13419 22269
rect 15929 22266 15995 22269
rect 11789 22264 15995 22266
rect 11789 22208 11794 22264
rect 11850 22208 13358 22264
rect 13414 22208 15934 22264
rect 15990 22208 15995 22264
rect 11789 22206 15995 22208
rect 11789 22203 11855 22206
rect 13353 22203 13419 22206
rect 15929 22203 15995 22206
rect 6269 22132 6335 22133
rect 6269 22130 6316 22132
rect 6224 22128 6316 22130
rect 6224 22072 6274 22128
rect 6224 22070 6316 22072
rect 6269 22068 6316 22070
rect 6380 22068 6386 22132
rect 7465 22130 7531 22133
rect 7465 22128 7850 22130
rect 7465 22072 7470 22128
rect 7526 22072 7850 22128
rect 7465 22070 7850 22072
rect 6269 22067 6335 22068
rect 7465 22067 7531 22070
rect 3233 21994 3299 21997
rect 5574 21994 5580 21996
rect 3233 21992 5580 21994
rect 3233 21936 3238 21992
rect 3294 21936 5580 21992
rect 3233 21934 5580 21936
rect 3233 21931 3299 21934
rect 5574 21932 5580 21934
rect 5644 21932 5650 21996
rect 5717 21994 5783 21997
rect 6269 21994 6335 21997
rect 5717 21992 6335 21994
rect 5717 21936 5722 21992
rect 5778 21936 6274 21992
rect 6330 21936 6335 21992
rect 5717 21934 6335 21936
rect 5717 21931 5783 21934
rect 6269 21931 6335 21934
rect 6545 21994 6611 21997
rect 6545 21992 7666 21994
rect 6545 21936 6550 21992
rect 6606 21936 7666 21992
rect 6545 21934 7666 21936
rect 6545 21931 6611 21934
rect 200 21858 800 21888
rect 1577 21858 1643 21861
rect 200 21856 1643 21858
rect 200 21800 1582 21856
rect 1638 21800 1643 21856
rect 200 21798 1643 21800
rect 200 21768 800 21798
rect 1577 21795 1643 21798
rect 5073 21858 5139 21861
rect 5717 21858 5783 21861
rect 5073 21856 5783 21858
rect 5073 21800 5078 21856
rect 5134 21800 5722 21856
rect 5778 21800 5783 21856
rect 5073 21798 5783 21800
rect 5073 21795 5139 21798
rect 5717 21795 5783 21798
rect 4429 21722 4495 21725
rect 5349 21722 5415 21725
rect 4429 21720 5415 21722
rect 4429 21664 4434 21720
rect 4490 21664 5354 21720
rect 5410 21664 5415 21720
rect 4429 21662 5415 21664
rect 7606 21722 7666 21934
rect 7790 21861 7850 22070
rect 9622 22068 9628 22132
rect 9692 22130 9698 22132
rect 16021 22130 16087 22133
rect 9692 22128 16087 22130
rect 9692 22072 16026 22128
rect 16082 22072 16087 22128
rect 9692 22070 16087 22072
rect 9692 22068 9698 22070
rect 16021 22067 16087 22070
rect 10777 21996 10843 21997
rect 10726 21994 10732 21996
rect 10686 21934 10732 21994
rect 10796 21992 10843 21996
rect 10838 21936 10843 21992
rect 10726 21932 10732 21934
rect 10796 21932 10843 21936
rect 10777 21931 10843 21932
rect 13261 21994 13327 21997
rect 14917 21994 14983 21997
rect 13261 21992 14983 21994
rect 13261 21936 13266 21992
rect 13322 21936 14922 21992
rect 14978 21936 14983 21992
rect 13261 21934 14983 21936
rect 13261 21931 13327 21934
rect 14917 21931 14983 21934
rect 7790 21856 7899 21861
rect 11053 21858 11119 21861
rect 7790 21800 7838 21856
rect 7894 21800 7899 21856
rect 7790 21798 7899 21800
rect 7833 21795 7899 21798
rect 9630 21856 11119 21858
rect 9630 21800 11058 21856
rect 11114 21800 11119 21856
rect 9630 21798 11119 21800
rect 9630 21722 9690 21798
rect 11053 21795 11119 21798
rect 11789 21858 11855 21861
rect 18321 21858 18387 21861
rect 11789 21856 18387 21858
rect 11789 21800 11794 21856
rect 11850 21800 18326 21856
rect 18382 21800 18387 21856
rect 11789 21798 18387 21800
rect 11789 21795 11855 21798
rect 18321 21795 18387 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 7606 21662 9690 21722
rect 10777 21722 10843 21725
rect 17677 21722 17743 21725
rect 10777 21720 17743 21722
rect 10777 21664 10782 21720
rect 10838 21664 17682 21720
rect 17738 21664 17743 21720
rect 10777 21662 17743 21664
rect 4429 21659 4495 21662
rect 5349 21659 5415 21662
rect 10777 21659 10843 21662
rect 17677 21659 17743 21662
rect 3877 21586 3943 21589
rect 4654 21586 4660 21588
rect 3877 21584 4660 21586
rect 3877 21528 3882 21584
rect 3938 21528 4660 21584
rect 3877 21526 4660 21528
rect 3877 21523 3943 21526
rect 4654 21524 4660 21526
rect 4724 21524 4730 21588
rect 10501 21586 10567 21589
rect 14181 21586 14247 21589
rect 10501 21584 14247 21586
rect 10501 21528 10506 21584
rect 10562 21528 14186 21584
rect 14242 21528 14247 21584
rect 10501 21526 14247 21528
rect 10501 21523 10567 21526
rect 14181 21523 14247 21526
rect 4245 21450 4311 21453
rect 6821 21450 6887 21453
rect 4245 21448 6887 21450
rect 4245 21392 4250 21448
rect 4306 21392 6826 21448
rect 6882 21392 6887 21448
rect 4245 21390 6887 21392
rect 4245 21387 4311 21390
rect 6821 21387 6887 21390
rect 19793 21450 19859 21453
rect 24393 21450 24459 21453
rect 19793 21448 24459 21450
rect 19793 21392 19798 21448
rect 19854 21392 24398 21448
rect 24454 21392 24459 21448
rect 19793 21390 24459 21392
rect 19793 21387 19859 21390
rect 24393 21387 24459 21390
rect 5441 21314 5507 21317
rect 5942 21314 5948 21316
rect 5441 21312 5948 21314
rect 5441 21256 5446 21312
rect 5502 21256 5948 21312
rect 5441 21254 5948 21256
rect 5441 21251 5507 21254
rect 5942 21252 5948 21254
rect 6012 21252 6018 21316
rect 9949 21314 10015 21317
rect 17493 21314 17559 21317
rect 9949 21312 17559 21314
rect 9949 21256 9954 21312
rect 10010 21256 17498 21312
rect 17554 21256 17559 21312
rect 9949 21254 17559 21256
rect 9949 21251 10015 21254
rect 17493 21251 17559 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 11513 21178 11579 21181
rect 7054 21176 11579 21178
rect 7054 21120 11518 21176
rect 11574 21120 11579 21176
rect 7054 21118 11579 21120
rect 6177 21042 6243 21045
rect 6310 21042 6316 21044
rect 6177 21040 6316 21042
rect 6177 20984 6182 21040
rect 6238 20984 6316 21040
rect 6177 20982 6316 20984
rect 6177 20979 6243 20982
rect 6310 20980 6316 20982
rect 6380 20980 6386 21044
rect 4521 20906 4587 20909
rect 6729 20906 6795 20909
rect 7054 20906 7114 21118
rect 11513 21115 11579 21118
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 10961 21042 11027 21045
rect 16573 21042 16639 21045
rect 10961 21040 16639 21042
rect 10961 20984 10966 21040
rect 11022 20984 16578 21040
rect 16634 20984 16639 21040
rect 10961 20982 16639 20984
rect 10961 20979 11027 20982
rect 16573 20979 16639 20982
rect 4521 20904 7114 20906
rect 4521 20848 4526 20904
rect 4582 20848 6734 20904
rect 6790 20848 7114 20904
rect 4521 20846 7114 20848
rect 8293 20906 8359 20909
rect 14222 20906 14228 20908
rect 8293 20904 14228 20906
rect 8293 20848 8298 20904
rect 8354 20848 14228 20904
rect 8293 20846 14228 20848
rect 4521 20843 4587 20846
rect 6729 20843 6795 20846
rect 8293 20843 8359 20846
rect 14222 20844 14228 20846
rect 14292 20844 14298 20908
rect 20161 20906 20227 20909
rect 15150 20904 20227 20906
rect 15150 20848 20166 20904
rect 20222 20848 20227 20904
rect 15150 20846 20227 20848
rect 3785 20770 3851 20773
rect 7005 20770 7071 20773
rect 3785 20768 7071 20770
rect 3785 20712 3790 20768
rect 3846 20712 7010 20768
rect 7066 20712 7071 20768
rect 3785 20710 7071 20712
rect 3785 20707 3851 20710
rect 7005 20707 7071 20710
rect 11053 20770 11119 20773
rect 15150 20770 15210 20846
rect 20161 20843 20227 20846
rect 11053 20768 15210 20770
rect 11053 20712 11058 20768
rect 11114 20712 15210 20768
rect 11053 20710 15210 20712
rect 15285 20770 15351 20773
rect 17718 20770 17724 20772
rect 15285 20768 17724 20770
rect 15285 20712 15290 20768
rect 15346 20712 17724 20768
rect 15285 20710 17724 20712
rect 11053 20707 11119 20710
rect 15285 20707 15351 20710
rect 17718 20708 17724 20710
rect 17788 20708 17794 20772
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 2589 20634 2655 20637
rect 2814 20634 2820 20636
rect 2589 20632 2820 20634
rect 2589 20576 2594 20632
rect 2650 20576 2820 20632
rect 2589 20574 2820 20576
rect 2589 20571 2655 20574
rect 2814 20572 2820 20574
rect 2884 20572 2890 20636
rect 3969 20634 4035 20637
rect 11421 20634 11487 20637
rect 3969 20632 11487 20634
rect 3969 20576 3974 20632
rect 4030 20576 11426 20632
rect 11482 20576 11487 20632
rect 3969 20574 11487 20576
rect 3969 20571 4035 20574
rect 11421 20571 11487 20574
rect 200 20498 800 20528
rect 2957 20498 3023 20501
rect 200 20496 3023 20498
rect 200 20440 2962 20496
rect 3018 20440 3023 20496
rect 200 20438 3023 20440
rect 200 20408 800 20438
rect 2957 20435 3023 20438
rect 3182 20436 3188 20500
rect 3252 20498 3258 20500
rect 12566 20498 12572 20500
rect 3252 20438 12572 20498
rect 3252 20436 3258 20438
rect 12566 20436 12572 20438
rect 12636 20436 12642 20500
rect 15009 20498 15075 20501
rect 15837 20498 15903 20501
rect 15009 20496 15903 20498
rect 15009 20440 15014 20496
rect 15070 20440 15842 20496
rect 15898 20440 15903 20496
rect 15009 20438 15903 20440
rect 15009 20435 15075 20438
rect 15837 20435 15903 20438
rect 37181 20498 37247 20501
rect 39200 20498 39800 20528
rect 37181 20496 39800 20498
rect 37181 20440 37186 20496
rect 37242 20440 39800 20496
rect 37181 20438 39800 20440
rect 37181 20435 37247 20438
rect 39200 20408 39800 20438
rect 5993 20362 6059 20365
rect 6453 20362 6519 20365
rect 13353 20362 13419 20365
rect 5993 20360 13419 20362
rect 5993 20304 5998 20360
rect 6054 20304 6458 20360
rect 6514 20304 13358 20360
rect 13414 20304 13419 20360
rect 5993 20302 13419 20304
rect 5993 20299 6059 20302
rect 6453 20299 6519 20302
rect 13353 20299 13419 20302
rect 14365 20362 14431 20365
rect 15653 20362 15719 20365
rect 14365 20360 15719 20362
rect 14365 20304 14370 20360
rect 14426 20304 15658 20360
rect 15714 20304 15719 20360
rect 14365 20302 15719 20304
rect 14365 20299 14431 20302
rect 15653 20299 15719 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 11421 20090 11487 20093
rect 17125 20090 17191 20093
rect 11421 20088 17191 20090
rect 11421 20032 11426 20088
rect 11482 20032 17130 20088
rect 17186 20032 17191 20088
rect 11421 20030 17191 20032
rect 11421 20027 11487 20030
rect 17125 20027 17191 20030
rect 9857 19954 9923 19957
rect 15653 19954 15719 19957
rect 9857 19952 15719 19954
rect 9857 19896 9862 19952
rect 9918 19896 15658 19952
rect 15714 19896 15719 19952
rect 9857 19894 15719 19896
rect 9857 19891 9923 19894
rect 15653 19891 15719 19894
rect 6177 19820 6243 19821
rect 6126 19818 6132 19820
rect 6050 19758 6132 19818
rect 6196 19818 6243 19820
rect 12934 19818 12940 19820
rect 6196 19816 12940 19818
rect 6238 19760 12940 19816
rect 6126 19756 6132 19758
rect 6196 19758 12940 19760
rect 6196 19756 6243 19758
rect 12934 19756 12940 19758
rect 13004 19756 13010 19820
rect 15469 19818 15535 19821
rect 18597 19818 18663 19821
rect 15469 19816 18663 19818
rect 15469 19760 15474 19816
rect 15530 19760 18602 19816
rect 18658 19760 18663 19816
rect 15469 19758 18663 19760
rect 6177 19755 6243 19756
rect 15469 19755 15535 19758
rect 18597 19755 18663 19758
rect 3601 19682 3667 19685
rect 10961 19682 11027 19685
rect 3601 19680 11027 19682
rect 3601 19624 3606 19680
rect 3662 19624 10966 19680
rect 11022 19624 11027 19680
rect 3601 19622 11027 19624
rect 3601 19619 3667 19622
rect 10961 19619 11027 19622
rect 11094 19620 11100 19684
rect 11164 19682 11170 19684
rect 11513 19682 11579 19685
rect 11646 19682 11652 19684
rect 11164 19680 11652 19682
rect 11164 19624 11518 19680
rect 11574 19624 11652 19680
rect 11164 19622 11652 19624
rect 11164 19620 11170 19622
rect 11513 19619 11579 19622
rect 11646 19620 11652 19622
rect 11716 19620 11722 19684
rect 12709 19682 12775 19685
rect 14457 19682 14523 19685
rect 12709 19680 14523 19682
rect 12709 19624 12714 19680
rect 12770 19624 14462 19680
rect 14518 19624 14523 19680
rect 12709 19622 14523 19624
rect 12709 19619 12775 19622
rect 14457 19619 14523 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 3693 19548 3759 19549
rect 1894 19484 1900 19548
rect 1964 19546 1970 19548
rect 1964 19486 2790 19546
rect 1964 19484 1970 19486
rect 2730 19274 2790 19486
rect 3693 19544 3740 19548
rect 3804 19546 3810 19548
rect 4337 19546 4403 19549
rect 7465 19546 7531 19549
rect 3693 19488 3698 19544
rect 3693 19484 3740 19488
rect 3804 19486 3850 19546
rect 4337 19544 7531 19546
rect 4337 19488 4342 19544
rect 4398 19488 7470 19544
rect 7526 19488 7531 19544
rect 4337 19486 7531 19488
rect 3804 19484 3810 19486
rect 3693 19483 3759 19484
rect 4337 19483 4403 19486
rect 7465 19483 7531 19486
rect 8385 19546 8451 19549
rect 15377 19546 15443 19549
rect 8385 19544 15443 19546
rect 8385 19488 8390 19544
rect 8446 19488 15382 19544
rect 15438 19488 15443 19544
rect 8385 19486 15443 19488
rect 8385 19483 8451 19486
rect 15377 19483 15443 19486
rect 7005 19412 7071 19413
rect 3918 19348 3924 19412
rect 3988 19410 3994 19412
rect 5022 19410 5028 19412
rect 3988 19350 5028 19410
rect 3988 19348 3994 19350
rect 5022 19348 5028 19350
rect 5092 19348 5098 19412
rect 7005 19408 7052 19412
rect 7116 19410 7122 19412
rect 9949 19410 10015 19413
rect 13997 19410 14063 19413
rect 7005 19352 7010 19408
rect 7005 19348 7052 19352
rect 7116 19350 7162 19410
rect 9949 19408 14063 19410
rect 9949 19352 9954 19408
rect 10010 19352 14002 19408
rect 14058 19352 14063 19408
rect 9949 19350 14063 19352
rect 7116 19348 7122 19350
rect 7005 19347 7071 19348
rect 9949 19347 10015 19350
rect 13997 19347 14063 19350
rect 9622 19274 9628 19276
rect 2730 19214 9628 19274
rect 9622 19212 9628 19214
rect 9692 19212 9698 19276
rect 10409 19274 10475 19277
rect 12433 19274 12499 19277
rect 10409 19272 12499 19274
rect 10409 19216 10414 19272
rect 10470 19216 12438 19272
rect 12494 19216 12499 19272
rect 10409 19214 12499 19216
rect 10409 19211 10475 19214
rect 12433 19211 12499 19214
rect 200 19138 800 19168
rect 7097 19138 7163 19141
rect 25129 19138 25195 19141
rect 25681 19138 25747 19141
rect 200 19078 2790 19138
rect 200 19048 800 19078
rect 2730 18866 2790 19078
rect 7097 19136 25747 19138
rect 7097 19080 7102 19136
rect 7158 19080 25134 19136
rect 25190 19080 25686 19136
rect 25742 19080 25747 19136
rect 7097 19078 25747 19080
rect 7097 19075 7163 19078
rect 25129 19075 25195 19078
rect 25681 19075 25747 19078
rect 38285 19138 38351 19141
rect 39200 19138 39800 19168
rect 38285 19136 39800 19138
rect 38285 19080 38290 19136
rect 38346 19080 39800 19136
rect 38285 19078 39800 19080
rect 38285 19075 38351 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 7281 19002 7347 19005
rect 11053 19002 11119 19005
rect 7281 19000 11119 19002
rect 7281 18944 7286 19000
rect 7342 18944 11058 19000
rect 11114 18944 11119 19000
rect 7281 18942 11119 18944
rect 7281 18939 7347 18942
rect 11053 18939 11119 18942
rect 5165 18866 5231 18869
rect 2730 18864 5231 18866
rect 2730 18808 5170 18864
rect 5226 18808 5231 18864
rect 2730 18806 5231 18808
rect 5165 18803 5231 18806
rect 6821 18866 6887 18869
rect 8845 18866 8911 18869
rect 6821 18864 8911 18866
rect 6821 18808 6826 18864
rect 6882 18808 8850 18864
rect 8906 18808 8911 18864
rect 6821 18806 8911 18808
rect 6821 18803 6887 18806
rect 8845 18803 8911 18806
rect 10225 18866 10291 18869
rect 10869 18866 10935 18869
rect 10225 18864 10935 18866
rect 10225 18808 10230 18864
rect 10286 18808 10874 18864
rect 10930 18808 10935 18864
rect 10225 18806 10935 18808
rect 10225 18803 10291 18806
rect 10869 18803 10935 18806
rect 11421 18866 11487 18869
rect 12065 18866 12131 18869
rect 12566 18866 12572 18868
rect 11421 18864 12572 18866
rect 11421 18808 11426 18864
rect 11482 18808 12070 18864
rect 12126 18808 12572 18864
rect 11421 18806 12572 18808
rect 11421 18803 11487 18806
rect 12065 18803 12131 18806
rect 12566 18804 12572 18806
rect 12636 18804 12642 18868
rect 8109 18730 8175 18733
rect 12157 18730 12223 18733
rect 8109 18728 12223 18730
rect 8109 18672 8114 18728
rect 8170 18672 12162 18728
rect 12218 18672 12223 18728
rect 8109 18670 12223 18672
rect 8109 18667 8175 18670
rect 12157 18667 12223 18670
rect 3325 18594 3391 18597
rect 6269 18594 6335 18597
rect 3325 18592 6335 18594
rect 3325 18536 3330 18592
rect 3386 18536 6274 18592
rect 6330 18536 6335 18592
rect 3325 18534 6335 18536
rect 3325 18531 3391 18534
rect 6269 18531 6335 18534
rect 6678 18532 6684 18596
rect 6748 18594 6754 18596
rect 7097 18594 7163 18597
rect 6748 18592 7163 18594
rect 6748 18536 7102 18592
rect 7158 18536 7163 18592
rect 6748 18534 7163 18536
rect 6748 18532 6754 18534
rect 7097 18531 7163 18534
rect 8937 18594 9003 18597
rect 11421 18594 11487 18597
rect 8937 18592 11487 18594
rect 8937 18536 8942 18592
rect 8998 18536 11426 18592
rect 11482 18536 11487 18592
rect 8937 18534 11487 18536
rect 8937 18531 9003 18534
rect 11421 18531 11487 18534
rect 11973 18594 12039 18597
rect 13445 18594 13511 18597
rect 11973 18592 13511 18594
rect 11973 18536 11978 18592
rect 12034 18536 13450 18592
rect 13506 18536 13511 18592
rect 11973 18534 13511 18536
rect 11973 18531 12039 18534
rect 13445 18531 13511 18534
rect 14038 18532 14044 18596
rect 14108 18594 14114 18596
rect 14181 18594 14247 18597
rect 14108 18592 14247 18594
rect 14108 18536 14186 18592
rect 14242 18536 14247 18592
rect 14108 18534 14247 18536
rect 14108 18532 14114 18534
rect 14181 18531 14247 18534
rect 19570 18528 19886 18529
rect 200 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 3233 18458 3299 18461
rect 200 18456 3299 18458
rect 200 18400 3238 18456
rect 3294 18400 3299 18456
rect 200 18398 3299 18400
rect 200 18368 800 18398
rect 3233 18395 3299 18398
rect 9857 18458 9923 18461
rect 12341 18458 12407 18461
rect 9857 18456 12407 18458
rect 9857 18400 9862 18456
rect 9918 18400 12346 18456
rect 12402 18400 12407 18456
rect 9857 18398 12407 18400
rect 9857 18395 9923 18398
rect 12341 18395 12407 18398
rect 13813 18458 13879 18461
rect 19241 18458 19307 18461
rect 13813 18456 19307 18458
rect 13813 18400 13818 18456
rect 13874 18400 19246 18456
rect 19302 18400 19307 18456
rect 13813 18398 19307 18400
rect 13813 18395 13879 18398
rect 19241 18395 19307 18398
rect 7005 18322 7071 18325
rect 7230 18322 7236 18324
rect 7005 18320 7236 18322
rect 7005 18264 7010 18320
rect 7066 18264 7236 18320
rect 7005 18262 7236 18264
rect 7005 18259 7071 18262
rect 7230 18260 7236 18262
rect 7300 18260 7306 18324
rect 12985 18322 13051 18325
rect 14549 18322 14615 18325
rect 12985 18320 14615 18322
rect 12985 18264 12990 18320
rect 13046 18264 14554 18320
rect 14610 18264 14615 18320
rect 12985 18262 14615 18264
rect 12985 18259 13051 18262
rect 14549 18259 14615 18262
rect 13445 18186 13511 18189
rect 15009 18186 15075 18189
rect 13445 18184 15075 18186
rect 13445 18128 13450 18184
rect 13506 18128 15014 18184
rect 15070 18128 15075 18184
rect 13445 18126 15075 18128
rect 13445 18123 13511 18126
rect 15009 18123 15075 18126
rect 5717 18052 5783 18053
rect 5717 18050 5764 18052
rect 5672 18048 5764 18050
rect 5672 17992 5722 18048
rect 5672 17990 5764 17992
rect 5717 17988 5764 17990
rect 5828 17988 5834 18052
rect 12065 18050 12131 18053
rect 16849 18050 16915 18053
rect 17350 18050 17356 18052
rect 12065 18048 17356 18050
rect 12065 17992 12070 18048
rect 12126 17992 16854 18048
rect 16910 17992 17356 18048
rect 12065 17990 17356 17992
rect 5717 17987 5783 17988
rect 12065 17987 12131 17990
rect 16849 17987 16915 17990
rect 17350 17988 17356 17990
rect 17420 17988 17426 18052
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 3325 17916 3391 17917
rect 3325 17912 3372 17916
rect 3436 17914 3442 17916
rect 10869 17914 10935 17917
rect 17861 17914 17927 17917
rect 3325 17856 3330 17912
rect 3325 17852 3372 17856
rect 3436 17854 3482 17914
rect 10869 17912 17927 17914
rect 10869 17856 10874 17912
rect 10930 17856 17866 17912
rect 17922 17856 17927 17912
rect 10869 17854 17927 17856
rect 3436 17852 3442 17854
rect 3325 17851 3391 17852
rect 10869 17851 10935 17854
rect 17861 17851 17927 17854
rect 3969 17778 4035 17781
rect 5441 17778 5507 17781
rect 3969 17776 5507 17778
rect 3969 17720 3974 17776
rect 4030 17720 5446 17776
rect 5502 17720 5507 17776
rect 3969 17718 5507 17720
rect 3969 17715 4035 17718
rect 5441 17715 5507 17718
rect 8937 17778 9003 17781
rect 9765 17778 9831 17781
rect 8937 17776 9831 17778
rect 8937 17720 8942 17776
rect 8998 17720 9770 17776
rect 9826 17720 9831 17776
rect 8937 17718 9831 17720
rect 8937 17715 9003 17718
rect 9765 17715 9831 17718
rect 11881 17778 11947 17781
rect 15285 17778 15351 17781
rect 11881 17776 15351 17778
rect 11881 17720 11886 17776
rect 11942 17720 15290 17776
rect 15346 17720 15351 17776
rect 11881 17718 15351 17720
rect 11881 17715 11947 17718
rect 15285 17715 15351 17718
rect 38193 17778 38259 17781
rect 39200 17778 39800 17808
rect 38193 17776 39800 17778
rect 38193 17720 38198 17776
rect 38254 17720 39800 17776
rect 38193 17718 39800 17720
rect 38193 17715 38259 17718
rect 39200 17688 39800 17718
rect 4521 17642 4587 17645
rect 6085 17642 6151 17645
rect 4521 17640 6151 17642
rect 4521 17584 4526 17640
rect 4582 17584 6090 17640
rect 6146 17584 6151 17640
rect 4521 17582 6151 17584
rect 4521 17579 4587 17582
rect 6085 17579 6151 17582
rect 3785 17506 3851 17509
rect 10225 17506 10291 17509
rect 3785 17504 10291 17506
rect 3785 17448 3790 17504
rect 3846 17448 10230 17504
rect 10286 17448 10291 17504
rect 3785 17446 10291 17448
rect 3785 17443 3851 17446
rect 10225 17443 10291 17446
rect 10869 17506 10935 17509
rect 13813 17506 13879 17509
rect 10869 17504 13879 17506
rect 10869 17448 10874 17504
rect 10930 17448 13818 17504
rect 13874 17448 13879 17504
rect 10869 17446 13879 17448
rect 10869 17443 10935 17446
rect 13813 17443 13879 17446
rect 15377 17506 15443 17509
rect 16246 17506 16252 17508
rect 15377 17504 16252 17506
rect 15377 17448 15382 17504
rect 15438 17448 16252 17504
rect 15377 17446 16252 17448
rect 15377 17443 15443 17446
rect 16246 17444 16252 17446
rect 16316 17444 16322 17508
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 1710 17308 1716 17372
rect 1780 17370 1786 17372
rect 1853 17370 1919 17373
rect 1780 17368 1919 17370
rect 1780 17312 1858 17368
rect 1914 17312 1919 17368
rect 1780 17310 1919 17312
rect 1780 17308 1786 17310
rect 1853 17307 1919 17310
rect 5993 17370 6059 17373
rect 6453 17370 6519 17373
rect 13629 17370 13695 17373
rect 5993 17368 13695 17370
rect 5993 17312 5998 17368
rect 6054 17312 6458 17368
rect 6514 17312 13634 17368
rect 13690 17312 13695 17368
rect 5993 17310 13695 17312
rect 5993 17307 6059 17310
rect 6453 17307 6519 17310
rect 13629 17307 13695 17310
rect 5441 17234 5507 17237
rect 13721 17234 13787 17237
rect 20161 17236 20227 17237
rect 20110 17234 20116 17236
rect 5441 17232 13787 17234
rect 5441 17176 5446 17232
rect 5502 17176 13726 17232
rect 13782 17176 13787 17232
rect 5441 17174 13787 17176
rect 20070 17174 20116 17234
rect 20180 17232 20227 17236
rect 20222 17176 20227 17232
rect 5441 17171 5507 17174
rect 13721 17171 13787 17174
rect 20110 17172 20116 17174
rect 20180 17172 20227 17176
rect 20161 17171 20227 17172
rect 200 17098 800 17128
rect 4889 17098 4955 17101
rect 200 17096 4955 17098
rect 200 17040 4894 17096
rect 4950 17040 4955 17096
rect 200 17038 4955 17040
rect 200 17008 800 17038
rect 4889 17035 4955 17038
rect 6729 17098 6795 17101
rect 23841 17098 23907 17101
rect 6729 17096 23907 17098
rect 6729 17040 6734 17096
rect 6790 17040 23846 17096
rect 23902 17040 23907 17096
rect 6729 17038 23907 17040
rect 6729 17035 6795 17038
rect 23841 17035 23907 17038
rect 3601 16962 3667 16965
rect 9397 16964 9463 16965
rect 3918 16962 3924 16964
rect 3601 16960 3924 16962
rect 3601 16904 3606 16960
rect 3662 16904 3924 16960
rect 3601 16902 3924 16904
rect 3601 16899 3667 16902
rect 3918 16900 3924 16902
rect 3988 16900 3994 16964
rect 9397 16960 9444 16964
rect 9508 16962 9514 16964
rect 10869 16962 10935 16965
rect 16573 16962 16639 16965
rect 9397 16904 9402 16960
rect 9397 16900 9444 16904
rect 9508 16902 9554 16962
rect 10869 16960 16639 16962
rect 10869 16904 10874 16960
rect 10930 16904 16578 16960
rect 16634 16904 16639 16960
rect 10869 16902 16639 16904
rect 9508 16900 9514 16902
rect 9397 16899 9463 16900
rect 10869 16899 10935 16902
rect 16573 16899 16639 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 9305 16826 9371 16829
rect 9581 16826 9647 16829
rect 9305 16824 9647 16826
rect 9305 16768 9310 16824
rect 9366 16768 9586 16824
rect 9642 16768 9647 16824
rect 9305 16766 9647 16768
rect 9305 16763 9371 16766
rect 9581 16763 9647 16766
rect 12341 16826 12407 16829
rect 16113 16826 16179 16829
rect 12341 16824 16179 16826
rect 12341 16768 12346 16824
rect 12402 16768 16118 16824
rect 16174 16768 16179 16824
rect 12341 16766 16179 16768
rect 12341 16763 12407 16766
rect 16113 16763 16179 16766
rect 9121 16690 9187 16693
rect 9305 16690 9371 16693
rect 10961 16692 11027 16693
rect 10910 16690 10916 16692
rect 9121 16688 9371 16690
rect 9121 16632 9126 16688
rect 9182 16632 9310 16688
rect 9366 16632 9371 16688
rect 9121 16630 9371 16632
rect 10870 16630 10916 16690
rect 10980 16688 11027 16692
rect 11022 16632 11027 16688
rect 9121 16627 9187 16630
rect 9305 16627 9371 16630
rect 10910 16628 10916 16630
rect 10980 16628 11027 16632
rect 10961 16627 11027 16628
rect 11605 16690 11671 16693
rect 13813 16690 13879 16693
rect 11605 16688 13879 16690
rect 11605 16632 11610 16688
rect 11666 16632 13818 16688
rect 13874 16632 13879 16688
rect 11605 16630 13879 16632
rect 11605 16627 11671 16630
rect 13813 16627 13879 16630
rect 7189 16556 7255 16557
rect 7189 16552 7236 16556
rect 7300 16554 7306 16556
rect 7649 16554 7715 16557
rect 9581 16554 9647 16557
rect 7189 16496 7194 16552
rect 7189 16492 7236 16496
rect 7300 16494 7346 16554
rect 7649 16552 9647 16554
rect 7649 16496 7654 16552
rect 7710 16496 9586 16552
rect 9642 16496 9647 16552
rect 7649 16494 9647 16496
rect 7300 16492 7306 16494
rect 7189 16491 7255 16492
rect 7649 16491 7715 16494
rect 9581 16491 9647 16494
rect 10501 16418 10567 16421
rect 14089 16418 14155 16421
rect 10501 16416 14155 16418
rect 10501 16360 10506 16416
rect 10562 16360 14094 16416
rect 14150 16360 14155 16416
rect 10501 16358 14155 16360
rect 10501 16355 10567 16358
rect 14089 16355 14155 16358
rect 38193 16418 38259 16421
rect 39200 16418 39800 16448
rect 38193 16416 39800 16418
rect 38193 16360 38198 16416
rect 38254 16360 39800 16416
rect 38193 16358 39800 16360
rect 38193 16355 38259 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 39200 16328 39800 16358
rect 19570 16287 19886 16288
rect 3785 16282 3851 16285
rect 6494 16282 6500 16284
rect 3785 16280 6500 16282
rect 3785 16224 3790 16280
rect 3846 16224 6500 16280
rect 3785 16222 6500 16224
rect 3785 16219 3851 16222
rect 6494 16220 6500 16222
rect 6564 16282 6570 16284
rect 7649 16282 7715 16285
rect 6564 16280 7715 16282
rect 6564 16224 7654 16280
rect 7710 16224 7715 16280
rect 6564 16222 7715 16224
rect 6564 16220 6570 16222
rect 7649 16219 7715 16222
rect 8150 16220 8156 16284
rect 8220 16282 8226 16284
rect 10409 16282 10475 16285
rect 8220 16280 10475 16282
rect 8220 16224 10414 16280
rect 10470 16224 10475 16280
rect 8220 16222 10475 16224
rect 8220 16220 8226 16222
rect 10409 16219 10475 16222
rect 13353 16282 13419 16285
rect 15285 16282 15351 16285
rect 13353 16280 15351 16282
rect 13353 16224 13358 16280
rect 13414 16224 15290 16280
rect 15346 16224 15351 16280
rect 13353 16222 15351 16224
rect 13353 16219 13419 16222
rect 15285 16219 15351 16222
rect 9765 16146 9831 16149
rect 11697 16146 11763 16149
rect 9765 16144 11763 16146
rect 9765 16088 9770 16144
rect 9826 16088 11702 16144
rect 11758 16088 11763 16144
rect 9765 16086 11763 16088
rect 9765 16083 9831 16086
rect 11697 16083 11763 16086
rect 12065 16146 12131 16149
rect 27613 16146 27679 16149
rect 12065 16144 27679 16146
rect 12065 16088 12070 16144
rect 12126 16088 27618 16144
rect 27674 16088 27679 16144
rect 12065 16086 27679 16088
rect 12065 16083 12131 16086
rect 27613 16083 27679 16086
rect 10961 15874 11027 15877
rect 13353 15874 13419 15877
rect 14273 15874 14339 15877
rect 10961 15872 14339 15874
rect 10961 15816 10966 15872
rect 11022 15816 13358 15872
rect 13414 15816 14278 15872
rect 14334 15816 14339 15872
rect 10961 15814 14339 15816
rect 10961 15811 11027 15814
rect 13353 15811 13419 15814
rect 14273 15811 14339 15814
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 2773 15738 2839 15741
rect 200 15736 2839 15738
rect 200 15680 2778 15736
rect 2834 15680 2839 15736
rect 200 15678 2839 15680
rect 200 15648 800 15678
rect 2773 15675 2839 15678
rect 11329 15738 11395 15741
rect 15561 15738 15627 15741
rect 11329 15736 15627 15738
rect 11329 15680 11334 15736
rect 11390 15680 15566 15736
rect 15622 15680 15627 15736
rect 11329 15678 15627 15680
rect 11329 15675 11395 15678
rect 15561 15675 15627 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 8109 15602 8175 15605
rect 12341 15602 12407 15605
rect 8109 15600 12407 15602
rect 8109 15544 8114 15600
rect 8170 15544 12346 15600
rect 12402 15544 12407 15600
rect 8109 15542 12407 15544
rect 8109 15539 8175 15542
rect 12341 15539 12407 15542
rect 12566 15540 12572 15604
rect 12636 15602 12642 15604
rect 13353 15602 13419 15605
rect 12636 15600 13419 15602
rect 12636 15544 13358 15600
rect 13414 15544 13419 15600
rect 12636 15542 13419 15544
rect 12636 15540 12642 15542
rect 13353 15539 13419 15542
rect 8753 15466 8819 15469
rect 21265 15466 21331 15469
rect 8753 15464 21331 15466
rect 8753 15408 8758 15464
rect 8814 15408 21270 15464
rect 21326 15408 21331 15464
rect 8753 15406 21331 15408
rect 8753 15403 8819 15406
rect 21265 15403 21331 15406
rect 3417 15330 3483 15333
rect 8385 15330 8451 15333
rect 9121 15330 9187 15333
rect 17125 15330 17191 15333
rect 3417 15328 9187 15330
rect 3417 15272 3422 15328
rect 3478 15272 8390 15328
rect 8446 15272 9126 15328
rect 9182 15272 9187 15328
rect 3417 15270 9187 15272
rect 3417 15267 3483 15270
rect 8385 15267 8451 15270
rect 9121 15267 9187 15270
rect 15150 15328 17191 15330
rect 15150 15272 17130 15328
rect 17186 15272 17191 15328
rect 15150 15270 17191 15272
rect 9305 15194 9371 15197
rect 12249 15194 12315 15197
rect 9305 15192 12315 15194
rect 9305 15136 9310 15192
rect 9366 15136 12254 15192
rect 12310 15136 12315 15192
rect 9305 15134 12315 15136
rect 9305 15131 9371 15134
rect 12249 15131 12315 15134
rect 12525 15194 12591 15197
rect 15150 15194 15210 15270
rect 17125 15267 17191 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 12525 15192 15210 15194
rect 12525 15136 12530 15192
rect 12586 15136 15210 15192
rect 12525 15134 15210 15136
rect 15469 15196 15535 15197
rect 15469 15192 15516 15196
rect 15580 15194 15586 15196
rect 15469 15136 15474 15192
rect 12525 15131 12591 15134
rect 15469 15132 15516 15136
rect 15580 15134 15626 15194
rect 15580 15132 15586 15134
rect 15469 15131 15535 15132
rect 200 15058 800 15088
rect 7097 15058 7163 15061
rect 200 15056 7163 15058
rect 200 15000 7102 15056
rect 7158 15000 7163 15056
rect 200 14998 7163 15000
rect 200 14968 800 14998
rect 7097 14995 7163 14998
rect 15009 15058 15075 15061
rect 17585 15058 17651 15061
rect 15009 15056 17651 15058
rect 15009 15000 15014 15056
rect 15070 15000 17590 15056
rect 17646 15000 17651 15056
rect 15009 14998 17651 15000
rect 15009 14995 15075 14998
rect 17585 14995 17651 14998
rect 3325 14922 3391 14925
rect 10726 14922 10732 14924
rect 3325 14920 10732 14922
rect 3325 14864 3330 14920
rect 3386 14864 10732 14920
rect 3325 14862 10732 14864
rect 3325 14859 3391 14862
rect 10726 14860 10732 14862
rect 10796 14922 10802 14924
rect 16113 14922 16179 14925
rect 10796 14920 16179 14922
rect 10796 14864 16118 14920
rect 16174 14864 16179 14920
rect 10796 14862 16179 14864
rect 10796 14860 10802 14862
rect 16113 14859 16179 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 11145 14650 11211 14653
rect 12065 14650 12131 14653
rect 11145 14648 12131 14650
rect 11145 14592 11150 14648
rect 11206 14592 12070 14648
rect 12126 14592 12131 14648
rect 11145 14590 12131 14592
rect 11145 14587 11211 14590
rect 12065 14587 12131 14590
rect 16246 14588 16252 14652
rect 16316 14650 16322 14652
rect 24669 14650 24735 14653
rect 16316 14648 24735 14650
rect 16316 14592 24674 14648
rect 24730 14592 24735 14648
rect 16316 14590 24735 14592
rect 16316 14588 16322 14590
rect 24669 14587 24735 14590
rect 8845 14514 8911 14517
rect 23197 14514 23263 14517
rect 8845 14512 23263 14514
rect 8845 14456 8850 14512
rect 8906 14456 23202 14512
rect 23258 14456 23263 14512
rect 8845 14454 23263 14456
rect 8845 14451 8911 14454
rect 23197 14451 23263 14454
rect 9489 14380 9555 14381
rect 9438 14316 9444 14380
rect 9508 14378 9555 14380
rect 10685 14378 10751 14381
rect 38193 14378 38259 14381
rect 39200 14378 39800 14408
rect 9508 14376 9600 14378
rect 9550 14320 9600 14376
rect 9508 14318 9600 14320
rect 10685 14376 11714 14378
rect 10685 14320 10690 14376
rect 10746 14320 11714 14376
rect 10685 14318 11714 14320
rect 9508 14316 9555 14318
rect 9489 14315 9555 14316
rect 10685 14315 10751 14318
rect 11654 14245 11714 14318
rect 38193 14376 39800 14378
rect 38193 14320 38198 14376
rect 38254 14320 39800 14376
rect 38193 14318 39800 14320
rect 38193 14315 38259 14318
rect 39200 14288 39800 14318
rect 11654 14240 11763 14245
rect 11654 14184 11702 14240
rect 11758 14184 11763 14240
rect 11654 14182 11763 14184
rect 11697 14179 11763 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 10041 14106 10107 14109
rect 18137 14106 18203 14109
rect 10041 14104 18203 14106
rect 10041 14048 10046 14104
rect 10102 14048 18142 14104
rect 18198 14048 18203 14104
rect 10041 14046 18203 14048
rect 10041 14043 10107 14046
rect 18137 14043 18203 14046
rect 8845 13834 8911 13837
rect 14038 13834 14044 13836
rect 8845 13832 14044 13834
rect 8845 13776 8850 13832
rect 8906 13776 14044 13832
rect 8845 13774 14044 13776
rect 8845 13771 8911 13774
rect 14038 13772 14044 13774
rect 14108 13772 14114 13836
rect 200 13698 800 13728
rect 2221 13698 2287 13701
rect 14273 13700 14339 13701
rect 200 13696 2287 13698
rect 200 13640 2226 13696
rect 2282 13640 2287 13696
rect 200 13638 2287 13640
rect 200 13608 800 13638
rect 2221 13635 2287 13638
rect 14222 13636 14228 13700
rect 14292 13698 14339 13700
rect 14292 13696 14384 13698
rect 14334 13640 14384 13696
rect 14292 13638 14384 13640
rect 14292 13636 14339 13638
rect 14273 13635 14339 13636
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 17953 13562 18019 13565
rect 18086 13562 18092 13564
rect 17953 13560 18092 13562
rect 17953 13504 17958 13560
rect 18014 13504 18092 13560
rect 17953 13502 18092 13504
rect 17953 13499 18019 13502
rect 18086 13500 18092 13502
rect 18156 13500 18162 13564
rect 5533 13426 5599 13429
rect 5901 13426 5967 13429
rect 15745 13426 15811 13429
rect 5533 13424 15811 13426
rect 5533 13368 5538 13424
rect 5594 13368 5906 13424
rect 5962 13368 15750 13424
rect 15806 13368 15811 13424
rect 5533 13366 15811 13368
rect 5533 13363 5599 13366
rect 5901 13363 5967 13366
rect 15745 13363 15811 13366
rect 5717 13290 5783 13293
rect 8293 13290 8359 13293
rect 5717 13288 8359 13290
rect 5717 13232 5722 13288
rect 5778 13232 8298 13288
rect 8354 13232 8359 13288
rect 5717 13230 8359 13232
rect 5717 13227 5783 13230
rect 8293 13227 8359 13230
rect 11421 13290 11487 13293
rect 17033 13290 17099 13293
rect 23565 13290 23631 13293
rect 11421 13288 17099 13290
rect 11421 13232 11426 13288
rect 11482 13232 17038 13288
rect 17094 13232 17099 13288
rect 11421 13230 17099 13232
rect 11421 13227 11487 13230
rect 17033 13227 17099 13230
rect 17174 13288 23631 13290
rect 17174 13232 23570 13288
rect 23626 13232 23631 13288
rect 17174 13230 23631 13232
rect 10910 13154 10916 13156
rect 9630 13094 10916 13154
rect 9630 13021 9690 13094
rect 10910 13092 10916 13094
rect 10980 13154 10986 13156
rect 17174 13154 17234 13230
rect 23565 13227 23631 13230
rect 10980 13094 17234 13154
rect 10980 13092 10986 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 9581 13016 9690 13021
rect 9581 12960 9586 13016
rect 9642 12960 9690 13016
rect 9581 12958 9690 12960
rect 10225 13018 10291 13021
rect 10593 13018 10659 13021
rect 14917 13018 14983 13021
rect 16113 13018 16179 13021
rect 10225 13016 16179 13018
rect 10225 12960 10230 13016
rect 10286 12960 10598 13016
rect 10654 12960 14922 13016
rect 14978 12960 16118 13016
rect 16174 12960 16179 13016
rect 10225 12958 16179 12960
rect 9581 12955 9647 12958
rect 10225 12955 10291 12958
rect 10593 12955 10659 12958
rect 14917 12955 14983 12958
rect 16113 12955 16179 12958
rect 38193 13018 38259 13021
rect 39200 13018 39800 13048
rect 38193 13016 39800 13018
rect 38193 12960 38198 13016
rect 38254 12960 39800 13016
rect 38193 12958 39800 12960
rect 38193 12955 38259 12958
rect 39200 12928 39800 12958
rect 4061 12882 4127 12885
rect 23381 12882 23447 12885
rect 4061 12880 23447 12882
rect 4061 12824 4066 12880
rect 4122 12824 23386 12880
rect 23442 12824 23447 12880
rect 4061 12822 23447 12824
rect 4061 12819 4127 12822
rect 23381 12819 23447 12822
rect 3325 12746 3391 12749
rect 8150 12746 8156 12748
rect 3325 12744 8156 12746
rect 3325 12688 3330 12744
rect 3386 12688 8156 12744
rect 3325 12686 8156 12688
rect 3325 12683 3391 12686
rect 8150 12684 8156 12686
rect 8220 12684 8226 12748
rect 11513 12746 11579 12749
rect 13169 12746 13235 12749
rect 11513 12744 13235 12746
rect 11513 12688 11518 12744
rect 11574 12688 13174 12744
rect 13230 12688 13235 12744
rect 11513 12686 13235 12688
rect 11513 12683 11579 12686
rect 13169 12683 13235 12686
rect 14273 12746 14339 12749
rect 15653 12746 15719 12749
rect 17033 12746 17099 12749
rect 14273 12744 17099 12746
rect 14273 12688 14278 12744
rect 14334 12688 15658 12744
rect 15714 12688 17038 12744
rect 17094 12688 17099 12744
rect 14273 12686 17099 12688
rect 14273 12683 14339 12686
rect 15653 12683 15719 12686
rect 17033 12683 17099 12686
rect 19609 12746 19675 12749
rect 20110 12746 20116 12748
rect 19609 12744 20116 12746
rect 19609 12688 19614 12744
rect 19670 12688 20116 12744
rect 19609 12686 20116 12688
rect 19609 12683 19675 12686
rect 20110 12684 20116 12686
rect 20180 12684 20186 12748
rect 6821 12610 6887 12613
rect 11145 12610 11211 12613
rect 13445 12610 13511 12613
rect 6821 12608 9138 12610
rect 6821 12552 6826 12608
rect 6882 12552 9138 12608
rect 6821 12550 9138 12552
rect 6821 12547 6887 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 7005 12474 7071 12477
rect 8569 12474 8635 12477
rect 7005 12472 8635 12474
rect 7005 12416 7010 12472
rect 7066 12416 8574 12472
rect 8630 12416 8635 12472
rect 7005 12414 8635 12416
rect 9078 12474 9138 12550
rect 11145 12608 13511 12610
rect 11145 12552 11150 12608
rect 11206 12552 13450 12608
rect 13506 12552 13511 12608
rect 11145 12550 13511 12552
rect 11145 12547 11211 12550
rect 13445 12547 13511 12550
rect 15101 12610 15167 12613
rect 21081 12610 21147 12613
rect 15101 12608 21147 12610
rect 15101 12552 15106 12608
rect 15162 12552 21086 12608
rect 21142 12552 21147 12608
rect 15101 12550 21147 12552
rect 15101 12547 15167 12550
rect 21081 12547 21147 12550
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 23289 12474 23355 12477
rect 9078 12472 23355 12474
rect 9078 12416 23294 12472
rect 23350 12416 23355 12472
rect 9078 12414 23355 12416
rect 7005 12411 7071 12414
rect 8569 12411 8635 12414
rect 23289 12411 23355 12414
rect 200 12338 800 12368
rect 3233 12338 3299 12341
rect 200 12336 3299 12338
rect 200 12280 3238 12336
rect 3294 12280 3299 12336
rect 200 12278 3299 12280
rect 200 12248 800 12278
rect 3233 12275 3299 12278
rect 7465 12338 7531 12341
rect 10225 12338 10291 12341
rect 7465 12336 10291 12338
rect 7465 12280 7470 12336
rect 7526 12280 10230 12336
rect 10286 12280 10291 12336
rect 7465 12278 10291 12280
rect 7465 12275 7531 12278
rect 10225 12275 10291 12278
rect 10409 12338 10475 12341
rect 12065 12338 12131 12341
rect 10409 12336 12131 12338
rect 10409 12280 10414 12336
rect 10470 12280 12070 12336
rect 12126 12280 12131 12336
rect 10409 12278 12131 12280
rect 10409 12275 10475 12278
rect 12065 12275 12131 12278
rect 16021 12338 16087 12341
rect 18137 12338 18203 12341
rect 16021 12336 18203 12338
rect 16021 12280 16026 12336
rect 16082 12280 18142 12336
rect 18198 12280 18203 12336
rect 16021 12278 18203 12280
rect 16021 12275 16087 12278
rect 18137 12275 18203 12278
rect 38285 12338 38351 12341
rect 39200 12338 39800 12368
rect 38285 12336 39800 12338
rect 38285 12280 38290 12336
rect 38346 12280 39800 12336
rect 38285 12278 39800 12280
rect 38285 12275 38351 12278
rect 39200 12248 39800 12278
rect 1117 12202 1183 12205
rect 4245 12202 4311 12205
rect 1117 12200 4311 12202
rect 1117 12144 1122 12200
rect 1178 12144 4250 12200
rect 4306 12144 4311 12200
rect 1117 12142 4311 12144
rect 1117 12139 1183 12142
rect 4245 12139 4311 12142
rect 5349 12202 5415 12205
rect 24853 12202 24919 12205
rect 5349 12200 24919 12202
rect 5349 12144 5354 12200
rect 5410 12144 24858 12200
rect 24914 12144 24919 12200
rect 5349 12142 24919 12144
rect 5349 12139 5415 12142
rect 24853 12139 24919 12142
rect 3969 12066 4035 12069
rect 11789 12066 11855 12069
rect 3969 12064 11855 12066
rect 3969 12008 3974 12064
rect 4030 12008 11794 12064
rect 11850 12008 11855 12064
rect 3969 12006 11855 12008
rect 3969 12003 4035 12006
rect 11789 12003 11855 12006
rect 14089 12066 14155 12069
rect 15193 12066 15259 12069
rect 14089 12064 15259 12066
rect 14089 12008 14094 12064
rect 14150 12008 15198 12064
rect 15254 12008 15259 12064
rect 14089 12006 15259 12008
rect 14089 12003 14155 12006
rect 15193 12003 15259 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 1853 11932 1919 11933
rect 1853 11930 1900 11932
rect 1772 11928 1900 11930
rect 1964 11930 1970 11932
rect 5901 11930 5967 11933
rect 1964 11928 5967 11930
rect 1772 11872 1858 11928
rect 1964 11872 5906 11928
rect 5962 11872 5967 11928
rect 1772 11870 1900 11872
rect 1853 11868 1900 11870
rect 1964 11870 5967 11872
rect 1964 11868 1970 11870
rect 1853 11867 1919 11868
rect 5901 11867 5967 11870
rect 11145 11930 11211 11933
rect 13629 11930 13695 11933
rect 11145 11928 13695 11930
rect 11145 11872 11150 11928
rect 11206 11872 13634 11928
rect 13690 11872 13695 11928
rect 11145 11870 13695 11872
rect 11145 11867 11211 11870
rect 13629 11867 13695 11870
rect 3918 11732 3924 11796
rect 3988 11794 3994 11796
rect 4521 11794 4587 11797
rect 23289 11794 23355 11797
rect 3988 11792 23355 11794
rect 3988 11736 4526 11792
rect 4582 11736 23294 11792
rect 23350 11736 23355 11792
rect 3988 11734 23355 11736
rect 3988 11732 3994 11734
rect 4521 11731 4587 11734
rect 23289 11731 23355 11734
rect 200 11658 800 11688
rect 2865 11658 2931 11661
rect 200 11656 2931 11658
rect 200 11600 2870 11656
rect 2926 11600 2931 11656
rect 200 11598 2931 11600
rect 200 11568 800 11598
rect 2865 11595 2931 11598
rect 9673 11658 9739 11661
rect 22553 11658 22619 11661
rect 9673 11656 22619 11658
rect 9673 11600 9678 11656
rect 9734 11600 22558 11656
rect 22614 11600 22619 11656
rect 9673 11598 22619 11600
rect 9673 11595 9739 11598
rect 22553 11595 22619 11598
rect 9949 11522 10015 11525
rect 16665 11522 16731 11525
rect 9949 11520 16731 11522
rect 9949 11464 9954 11520
rect 10010 11464 16670 11520
rect 16726 11464 16731 11520
rect 9949 11462 16731 11464
rect 9949 11459 10015 11462
rect 16665 11459 16731 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 7557 11386 7623 11389
rect 9305 11386 9371 11389
rect 7557 11384 9371 11386
rect 7557 11328 7562 11384
rect 7618 11328 9310 11384
rect 9366 11328 9371 11384
rect 7557 11326 9371 11328
rect 7557 11323 7623 11326
rect 9305 11323 9371 11326
rect 15469 11386 15535 11389
rect 18045 11386 18111 11389
rect 15469 11384 18111 11386
rect 15469 11328 15474 11384
rect 15530 11328 18050 11384
rect 18106 11328 18111 11384
rect 15469 11326 18111 11328
rect 15469 11323 15535 11326
rect 18045 11323 18111 11326
rect 11646 11188 11652 11252
rect 11716 11250 11722 11252
rect 15142 11250 15148 11252
rect 11716 11190 15148 11250
rect 11716 11188 11722 11190
rect 15142 11188 15148 11190
rect 15212 11250 15218 11252
rect 17217 11250 17283 11253
rect 15212 11248 17283 11250
rect 15212 11192 17222 11248
rect 17278 11192 17283 11248
rect 15212 11190 17283 11192
rect 15212 11188 15218 11190
rect 17217 11187 17283 11190
rect 10726 11052 10732 11116
rect 10796 11114 10802 11116
rect 11237 11114 11303 11117
rect 10796 11112 11303 11114
rect 10796 11056 11242 11112
rect 11298 11056 11303 11112
rect 10796 11054 11303 11056
rect 10796 11052 10802 11054
rect 11237 11051 11303 11054
rect 13670 11052 13676 11116
rect 13740 11114 13746 11116
rect 19977 11114 20043 11117
rect 13740 11112 20043 11114
rect 13740 11056 19982 11112
rect 20038 11056 20043 11112
rect 13740 11054 20043 11056
rect 13740 11052 13746 11054
rect 19977 11051 20043 11054
rect 21909 11114 21975 11117
rect 27337 11114 27403 11117
rect 21909 11112 27403 11114
rect 21909 11056 21914 11112
rect 21970 11056 27342 11112
rect 27398 11056 27403 11112
rect 21909 11054 27403 11056
rect 21909 11051 21975 11054
rect 27337 11051 27403 11054
rect 10593 10978 10659 10981
rect 13077 10978 13143 10981
rect 18689 10978 18755 10981
rect 10593 10976 18755 10978
rect 10593 10920 10598 10976
rect 10654 10920 13082 10976
rect 13138 10920 18694 10976
rect 18750 10920 18755 10976
rect 10593 10918 18755 10920
rect 10593 10915 10659 10918
rect 13077 10915 13143 10918
rect 18689 10915 18755 10918
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 2313 10842 2379 10845
rect 2446 10842 2452 10844
rect 2313 10840 2452 10842
rect 2313 10784 2318 10840
rect 2374 10784 2452 10840
rect 2313 10782 2452 10784
rect 2313 10779 2379 10782
rect 2446 10780 2452 10782
rect 2516 10780 2522 10844
rect 11329 10842 11395 10845
rect 13813 10842 13879 10845
rect 11329 10840 13879 10842
rect 11329 10784 11334 10840
rect 11390 10784 13818 10840
rect 13874 10784 13879 10840
rect 11329 10782 13879 10784
rect 11329 10779 11395 10782
rect 13813 10779 13879 10782
rect 19977 10842 20043 10845
rect 24117 10842 24183 10845
rect 19977 10840 24183 10842
rect 19977 10784 19982 10840
rect 20038 10784 24122 10840
rect 24178 10784 24183 10840
rect 19977 10782 24183 10784
rect 19977 10779 20043 10782
rect 24117 10779 24183 10782
rect 6821 10706 6887 10709
rect 17033 10706 17099 10709
rect 6821 10704 17099 10706
rect 6821 10648 6826 10704
rect 6882 10648 17038 10704
rect 17094 10648 17099 10704
rect 6821 10646 17099 10648
rect 6821 10643 6887 10646
rect 17033 10643 17099 10646
rect 19333 10706 19399 10709
rect 21541 10706 21607 10709
rect 19333 10704 21607 10706
rect 19333 10648 19338 10704
rect 19394 10648 21546 10704
rect 21602 10648 21607 10704
rect 19333 10646 21607 10648
rect 19333 10643 19399 10646
rect 21541 10643 21607 10646
rect 3601 10570 3667 10573
rect 23289 10570 23355 10573
rect 3601 10568 23355 10570
rect 3601 10512 3606 10568
rect 3662 10512 23294 10568
rect 23350 10512 23355 10568
rect 3601 10510 23355 10512
rect 3601 10507 3667 10510
rect 23289 10507 23355 10510
rect 19701 10434 19767 10437
rect 20253 10434 20319 10437
rect 19701 10432 20319 10434
rect 19701 10376 19706 10432
rect 19762 10376 20258 10432
rect 20314 10376 20319 10432
rect 19701 10374 20319 10376
rect 19701 10371 19767 10374
rect 20253 10371 20319 10374
rect 20989 10434 21055 10437
rect 22093 10434 22159 10437
rect 20989 10432 22159 10434
rect 20989 10376 20994 10432
rect 21050 10376 22098 10432
rect 22154 10376 22159 10432
rect 20989 10374 22159 10376
rect 20989 10371 21055 10374
rect 22093 10371 22159 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 2773 10298 2839 10301
rect 200 10296 2839 10298
rect 200 10240 2778 10296
rect 2834 10240 2839 10296
rect 200 10238 2839 10240
rect 200 10208 800 10238
rect 2773 10235 2839 10238
rect 17718 10236 17724 10300
rect 17788 10298 17794 10300
rect 23657 10298 23723 10301
rect 17788 10296 23723 10298
rect 17788 10240 23662 10296
rect 23718 10240 23723 10296
rect 17788 10238 23723 10240
rect 17788 10236 17794 10238
rect 23657 10235 23723 10238
rect 7833 10162 7899 10165
rect 8477 10162 8543 10165
rect 7833 10160 8543 10162
rect 7833 10104 7838 10160
rect 7894 10104 8482 10160
rect 8538 10104 8543 10160
rect 7833 10102 8543 10104
rect 7833 10099 7899 10102
rect 8477 10099 8543 10102
rect 11881 10162 11947 10165
rect 14273 10162 14339 10165
rect 11881 10160 14339 10162
rect 11881 10104 11886 10160
rect 11942 10104 14278 10160
rect 14334 10104 14339 10160
rect 11881 10102 14339 10104
rect 11881 10099 11947 10102
rect 14273 10099 14339 10102
rect 16573 10162 16639 10165
rect 25037 10162 25103 10165
rect 16573 10160 25103 10162
rect 16573 10104 16578 10160
rect 16634 10104 25042 10160
rect 25098 10104 25103 10160
rect 16573 10102 25103 10104
rect 16573 10099 16639 10102
rect 25037 10099 25103 10102
rect 11605 10026 11671 10029
rect 12157 10026 12223 10029
rect 21265 10026 21331 10029
rect 11605 10024 21331 10026
rect 11605 9968 11610 10024
rect 11666 9968 12162 10024
rect 12218 9968 21270 10024
rect 21326 9968 21331 10024
rect 11605 9966 21331 9968
rect 11605 9963 11671 9966
rect 12157 9963 12223 9966
rect 21265 9963 21331 9966
rect 21817 10026 21883 10029
rect 23841 10026 23907 10029
rect 21817 10024 23907 10026
rect 21817 9968 21822 10024
rect 21878 9968 23846 10024
rect 23902 9968 23907 10024
rect 21817 9966 23907 9968
rect 21817 9963 21883 9966
rect 23841 9963 23907 9966
rect 9673 9890 9739 9893
rect 18965 9890 19031 9893
rect 9673 9888 19031 9890
rect 9673 9832 9678 9888
rect 9734 9832 18970 9888
rect 19026 9832 19031 9888
rect 9673 9830 19031 9832
rect 9673 9827 9739 9830
rect 18965 9827 19031 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 5441 9754 5507 9757
rect 7046 9754 7052 9756
rect 5441 9752 7052 9754
rect 5441 9696 5446 9752
rect 5502 9696 7052 9752
rect 5441 9694 7052 9696
rect 5441 9691 5507 9694
rect 7046 9692 7052 9694
rect 7116 9692 7122 9756
rect 19977 9754 20043 9757
rect 22829 9754 22895 9757
rect 19977 9752 22895 9754
rect 19977 9696 19982 9752
rect 20038 9696 22834 9752
rect 22890 9696 22895 9752
rect 19977 9694 22895 9696
rect 19977 9691 20043 9694
rect 22829 9691 22895 9694
rect 9581 9618 9647 9621
rect 24393 9618 24459 9621
rect 9581 9616 24459 9618
rect 9581 9560 9586 9616
rect 9642 9560 24398 9616
rect 24454 9560 24459 9616
rect 9581 9558 24459 9560
rect 9581 9555 9647 9558
rect 24393 9555 24459 9558
rect 37181 9618 37247 9621
rect 39200 9618 39800 9648
rect 37181 9616 39800 9618
rect 37181 9560 37186 9616
rect 37242 9560 39800 9616
rect 37181 9558 39800 9560
rect 37181 9555 37247 9558
rect 39200 9528 39800 9558
rect 5022 9420 5028 9484
rect 5092 9482 5098 9484
rect 6545 9482 6611 9485
rect 5092 9480 6611 9482
rect 5092 9424 6550 9480
rect 6606 9424 6611 9480
rect 5092 9422 6611 9424
rect 5092 9420 5098 9422
rect 6545 9419 6611 9422
rect 11513 9482 11579 9485
rect 15326 9482 15332 9484
rect 11513 9480 15332 9482
rect 11513 9424 11518 9480
rect 11574 9424 15332 9480
rect 11513 9422 15332 9424
rect 11513 9419 11579 9422
rect 15326 9420 15332 9422
rect 15396 9482 15402 9484
rect 15929 9482 15995 9485
rect 15396 9480 15995 9482
rect 15396 9424 15934 9480
rect 15990 9424 15995 9480
rect 15396 9422 15995 9424
rect 15396 9420 15402 9422
rect 15929 9419 15995 9422
rect 19374 9420 19380 9484
rect 19444 9482 19450 9484
rect 23841 9482 23907 9485
rect 19444 9480 23907 9482
rect 19444 9424 23846 9480
rect 23902 9424 23907 9480
rect 19444 9422 23907 9424
rect 19444 9420 19450 9422
rect 23841 9419 23907 9422
rect 10869 9346 10935 9349
rect 23381 9346 23447 9349
rect 10869 9344 23447 9346
rect 10869 9288 10874 9344
rect 10930 9288 23386 9344
rect 23442 9288 23447 9344
rect 10869 9286 23447 9288
rect 10869 9283 10935 9286
rect 23381 9283 23447 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 2589 9212 2655 9213
rect 2589 9210 2636 9212
rect 2544 9208 2636 9210
rect 2544 9152 2594 9208
rect 2544 9150 2636 9152
rect 2589 9148 2636 9150
rect 2700 9148 2706 9212
rect 11789 9210 11855 9213
rect 12525 9210 12591 9213
rect 11789 9208 12591 9210
rect 11789 9152 11794 9208
rect 11850 9152 12530 9208
rect 12586 9152 12591 9208
rect 11789 9150 12591 9152
rect 2589 9147 2655 9148
rect 11789 9147 11855 9150
rect 12525 9147 12591 9150
rect 15745 9210 15811 9213
rect 23105 9210 23171 9213
rect 15745 9208 23171 9210
rect 15745 9152 15750 9208
rect 15806 9152 23110 9208
rect 23166 9152 23171 9208
rect 15745 9150 23171 9152
rect 15745 9147 15811 9150
rect 23105 9147 23171 9150
rect 3233 9074 3299 9077
rect 4061 9074 4127 9077
rect 25221 9074 25287 9077
rect 3233 9072 25287 9074
rect 3233 9016 3238 9072
rect 3294 9016 4066 9072
rect 4122 9016 25226 9072
rect 25282 9016 25287 9072
rect 3233 9014 25287 9016
rect 3233 9011 3299 9014
rect 4061 9011 4127 9014
rect 25221 9011 25287 9014
rect 200 8938 800 8968
rect 1761 8938 1827 8941
rect 200 8936 1827 8938
rect 200 8880 1766 8936
rect 1822 8880 1827 8936
rect 200 8878 1827 8880
rect 200 8848 800 8878
rect 1761 8875 1827 8878
rect 6729 8938 6795 8941
rect 10777 8938 10843 8941
rect 6729 8936 10843 8938
rect 6729 8880 6734 8936
rect 6790 8880 10782 8936
rect 10838 8880 10843 8936
rect 6729 8878 10843 8880
rect 6729 8875 6795 8878
rect 10777 8875 10843 8878
rect 11513 8938 11579 8941
rect 15009 8938 15075 8941
rect 11513 8936 15075 8938
rect 11513 8880 11518 8936
rect 11574 8880 15014 8936
rect 15070 8880 15075 8936
rect 11513 8878 15075 8880
rect 11513 8875 11579 8878
rect 15009 8875 15075 8878
rect 17769 8938 17835 8941
rect 19333 8938 19399 8941
rect 20294 8938 20300 8940
rect 17769 8936 20300 8938
rect 17769 8880 17774 8936
rect 17830 8880 19338 8936
rect 19394 8880 20300 8936
rect 17769 8878 20300 8880
rect 17769 8875 17835 8878
rect 19333 8875 19399 8878
rect 20294 8876 20300 8878
rect 20364 8876 20370 8940
rect 13261 8802 13327 8805
rect 14181 8802 14247 8805
rect 13261 8800 14247 8802
rect 13261 8744 13266 8800
rect 13322 8744 14186 8800
rect 14242 8744 14247 8800
rect 13261 8742 14247 8744
rect 13261 8739 13327 8742
rect 14181 8739 14247 8742
rect 18137 8802 18203 8805
rect 18873 8802 18939 8805
rect 18137 8800 18939 8802
rect 18137 8744 18142 8800
rect 18198 8744 18878 8800
rect 18934 8744 18939 8800
rect 18137 8742 18939 8744
rect 18137 8739 18203 8742
rect 18873 8739 18939 8742
rect 19333 8804 19399 8805
rect 20161 8804 20227 8805
rect 19333 8800 19380 8804
rect 19444 8802 19450 8804
rect 20110 8802 20116 8804
rect 19333 8744 19338 8800
rect 19333 8740 19380 8744
rect 19444 8742 19490 8802
rect 20070 8742 20116 8802
rect 20180 8800 20227 8804
rect 20222 8744 20227 8800
rect 19444 8740 19450 8742
rect 20110 8740 20116 8742
rect 20180 8740 20227 8744
rect 19333 8739 19399 8740
rect 20161 8739 20227 8740
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 10409 8666 10475 8669
rect 14089 8666 14155 8669
rect 10409 8664 14155 8666
rect 10409 8608 10414 8664
rect 10470 8608 14094 8664
rect 14150 8608 14155 8664
rect 10409 8606 14155 8608
rect 10409 8603 10475 8606
rect 14089 8603 14155 8606
rect 17309 8666 17375 8669
rect 18689 8666 18755 8669
rect 19057 8666 19123 8669
rect 17309 8664 19123 8666
rect 17309 8608 17314 8664
rect 17370 8608 18694 8664
rect 18750 8608 19062 8664
rect 19118 8608 19123 8664
rect 17309 8606 19123 8608
rect 17309 8603 17375 8606
rect 18689 8603 18755 8606
rect 19057 8603 19123 8606
rect 19977 8666 20043 8669
rect 25313 8666 25379 8669
rect 19977 8664 25379 8666
rect 19977 8608 19982 8664
rect 20038 8608 25318 8664
rect 25374 8608 25379 8664
rect 19977 8606 25379 8608
rect 19977 8603 20043 8606
rect 25313 8603 25379 8606
rect 22001 8530 22067 8533
rect 12390 8528 22067 8530
rect 12390 8472 22006 8528
rect 22062 8472 22067 8528
rect 12390 8470 22067 8472
rect 9213 8394 9279 8397
rect 12390 8394 12450 8470
rect 22001 8467 22067 8470
rect 9213 8392 12450 8394
rect 9213 8336 9218 8392
rect 9274 8336 12450 8392
rect 9213 8334 12450 8336
rect 9213 8331 9279 8334
rect 12934 8332 12940 8396
rect 13004 8394 13010 8396
rect 17585 8394 17651 8397
rect 13004 8392 17651 8394
rect 13004 8336 17590 8392
rect 17646 8336 17651 8392
rect 13004 8334 17651 8336
rect 13004 8332 13010 8334
rect 17585 8331 17651 8334
rect 19374 8332 19380 8396
rect 19444 8394 19450 8396
rect 20253 8394 20319 8397
rect 21725 8394 21791 8397
rect 19444 8392 21791 8394
rect 19444 8336 20258 8392
rect 20314 8336 21730 8392
rect 21786 8336 21791 8392
rect 19444 8334 21791 8336
rect 19444 8332 19450 8334
rect 20253 8331 20319 8334
rect 21725 8331 21791 8334
rect 8334 8196 8340 8260
rect 8404 8258 8410 8260
rect 8569 8258 8635 8261
rect 8404 8256 8635 8258
rect 8404 8200 8574 8256
rect 8630 8200 8635 8256
rect 8404 8198 8635 8200
rect 8404 8196 8410 8198
rect 8569 8195 8635 8198
rect 9673 8258 9739 8261
rect 12157 8258 12223 8261
rect 9673 8256 12223 8258
rect 9673 8200 9678 8256
rect 9734 8200 12162 8256
rect 12218 8200 12223 8256
rect 9673 8198 12223 8200
rect 9673 8195 9739 8198
rect 12157 8195 12223 8198
rect 17125 8258 17191 8261
rect 31385 8258 31451 8261
rect 17125 8256 31451 8258
rect 17125 8200 17130 8256
rect 17186 8200 31390 8256
rect 31446 8200 31451 8256
rect 17125 8198 31451 8200
rect 17125 8195 17191 8198
rect 31385 8195 31451 8198
rect 38285 8258 38351 8261
rect 39200 8258 39800 8288
rect 38285 8256 39800 8258
rect 38285 8200 38290 8256
rect 38346 8200 39800 8256
rect 38285 8198 39800 8200
rect 38285 8195 38351 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 10961 8122 11027 8125
rect 14549 8122 14615 8125
rect 10961 8120 14615 8122
rect 10961 8064 10966 8120
rect 11022 8064 14554 8120
rect 14610 8064 14615 8120
rect 10961 8062 14615 8064
rect 10961 8059 11027 8062
rect 14549 8059 14615 8062
rect 16573 8122 16639 8125
rect 22461 8122 22527 8125
rect 16573 8120 22527 8122
rect 16573 8064 16578 8120
rect 16634 8064 22466 8120
rect 22522 8064 22527 8120
rect 16573 8062 22527 8064
rect 16573 8059 16639 8062
rect 22461 8059 22527 8062
rect 2865 7986 2931 7989
rect 25221 7986 25287 7989
rect 2865 7984 25287 7986
rect 2865 7928 2870 7984
rect 2926 7928 25226 7984
rect 25282 7928 25287 7984
rect 2865 7926 25287 7928
rect 2865 7923 2931 7926
rect 25221 7923 25287 7926
rect 10409 7850 10475 7853
rect 13997 7850 14063 7853
rect 19885 7850 19951 7853
rect 10409 7848 19951 7850
rect 10409 7792 10414 7848
rect 10470 7792 14002 7848
rect 14058 7792 19890 7848
rect 19946 7792 19951 7848
rect 10409 7790 19951 7792
rect 10409 7787 10475 7790
rect 13997 7787 14063 7790
rect 19885 7787 19951 7790
rect 20069 7850 20135 7853
rect 22369 7850 22435 7853
rect 20069 7848 22435 7850
rect 20069 7792 20074 7848
rect 20130 7792 22374 7848
rect 22430 7792 22435 7848
rect 20069 7790 22435 7792
rect 20069 7787 20135 7790
rect 22369 7787 22435 7790
rect 11145 7714 11211 7717
rect 12065 7714 12131 7717
rect 17953 7714 18019 7717
rect 11145 7712 11346 7714
rect 11145 7656 11150 7712
rect 11206 7656 11346 7712
rect 11145 7654 11346 7656
rect 11145 7651 11211 7654
rect 200 7578 800 7608
rect 1577 7578 1643 7581
rect 200 7576 1643 7578
rect 200 7520 1582 7576
rect 1638 7520 1643 7576
rect 200 7518 1643 7520
rect 200 7488 800 7518
rect 1577 7515 1643 7518
rect 4797 7578 4863 7581
rect 11145 7578 11211 7581
rect 4797 7576 11211 7578
rect 4797 7520 4802 7576
rect 4858 7520 11150 7576
rect 11206 7520 11211 7576
rect 4797 7518 11211 7520
rect 11286 7578 11346 7654
rect 12065 7712 18019 7714
rect 12065 7656 12070 7712
rect 12126 7656 17958 7712
rect 18014 7656 18019 7712
rect 12065 7654 18019 7656
rect 12065 7651 12131 7654
rect 17953 7651 18019 7654
rect 19977 7714 20043 7717
rect 20437 7714 20503 7717
rect 19977 7712 20503 7714
rect 19977 7656 19982 7712
rect 20038 7656 20442 7712
rect 20498 7656 20503 7712
rect 19977 7654 20503 7656
rect 19977 7651 20043 7654
rect 20437 7651 20503 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 15469 7578 15535 7581
rect 11286 7576 15535 7578
rect 11286 7520 15474 7576
rect 15530 7520 15535 7576
rect 11286 7518 15535 7520
rect 4797 7515 4863 7518
rect 11145 7515 11211 7518
rect 15469 7515 15535 7518
rect 17677 7580 17743 7581
rect 17677 7576 17724 7580
rect 17788 7578 17794 7580
rect 23841 7578 23907 7581
rect 17677 7520 17682 7576
rect 17677 7516 17724 7520
rect 17788 7518 17834 7578
rect 20118 7576 23907 7578
rect 20118 7520 23846 7576
rect 23902 7520 23907 7576
rect 20118 7518 23907 7520
rect 17788 7516 17794 7518
rect 17677 7515 17743 7516
rect 10961 7442 11027 7445
rect 20118 7442 20178 7518
rect 23841 7515 23907 7518
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 10961 7440 20178 7442
rect 10961 7384 10966 7440
rect 11022 7384 20178 7440
rect 10961 7382 20178 7384
rect 20345 7442 20411 7445
rect 22921 7442 22987 7445
rect 20345 7440 22987 7442
rect 20345 7384 20350 7440
rect 20406 7384 22926 7440
rect 22982 7384 22987 7440
rect 20345 7382 22987 7384
rect 10961 7379 11027 7382
rect 20345 7379 20411 7382
rect 22921 7379 22987 7382
rect 6545 7306 6611 7309
rect 8845 7306 8911 7309
rect 6545 7304 8911 7306
rect 6545 7248 6550 7304
rect 6606 7248 8850 7304
rect 8906 7248 8911 7304
rect 6545 7246 8911 7248
rect 6545 7243 6611 7246
rect 8845 7243 8911 7246
rect 11053 7306 11119 7309
rect 24853 7306 24919 7309
rect 11053 7304 24919 7306
rect 11053 7248 11058 7304
rect 11114 7248 24858 7304
rect 24914 7248 24919 7304
rect 11053 7246 24919 7248
rect 11053 7243 11119 7246
rect 24853 7243 24919 7246
rect 7649 7170 7715 7173
rect 8753 7170 8819 7173
rect 7649 7168 8819 7170
rect 7649 7112 7654 7168
rect 7710 7112 8758 7168
rect 8814 7112 8819 7168
rect 7649 7110 8819 7112
rect 7649 7107 7715 7110
rect 8753 7107 8819 7110
rect 13486 7108 13492 7172
rect 13556 7170 13562 7172
rect 24853 7170 24919 7173
rect 13556 7168 24919 7170
rect 13556 7112 24858 7168
rect 24914 7112 24919 7168
rect 13556 7110 24919 7112
rect 13556 7108 13562 7110
rect 24853 7107 24919 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 9581 7034 9647 7037
rect 4846 7032 9647 7034
rect 4846 6976 9586 7032
rect 9642 6976 9647 7032
rect 4846 6974 9647 6976
rect 200 6898 800 6928
rect 4846 6898 4906 6974
rect 9581 6971 9647 6974
rect 16573 7034 16639 7037
rect 17350 7034 17356 7036
rect 16573 7032 17356 7034
rect 16573 6976 16578 7032
rect 16634 6976 17356 7032
rect 16573 6974 17356 6976
rect 16573 6971 16639 6974
rect 17350 6972 17356 6974
rect 17420 7034 17426 7036
rect 22001 7034 22067 7037
rect 17420 7032 22067 7034
rect 17420 6976 22006 7032
rect 22062 6976 22067 7032
rect 17420 6974 22067 6976
rect 17420 6972 17426 6974
rect 22001 6971 22067 6974
rect 200 6838 4906 6898
rect 6177 6898 6243 6901
rect 8569 6898 8635 6901
rect 6177 6896 8635 6898
rect 6177 6840 6182 6896
rect 6238 6840 8574 6896
rect 8630 6840 8635 6896
rect 6177 6838 8635 6840
rect 200 6808 800 6838
rect 6177 6835 6243 6838
rect 8569 6835 8635 6838
rect 9029 6898 9095 6901
rect 14641 6898 14707 6901
rect 9029 6896 14707 6898
rect 9029 6840 9034 6896
rect 9090 6840 14646 6896
rect 14702 6840 14707 6896
rect 9029 6838 14707 6840
rect 9029 6835 9095 6838
rect 14641 6835 14707 6838
rect 16757 6898 16823 6901
rect 26049 6898 26115 6901
rect 16757 6896 26115 6898
rect 16757 6840 16762 6896
rect 16818 6840 26054 6896
rect 26110 6840 26115 6896
rect 16757 6838 26115 6840
rect 16757 6835 16823 6838
rect 26049 6835 26115 6838
rect 6310 6700 6316 6764
rect 6380 6762 6386 6764
rect 9397 6762 9463 6765
rect 16113 6762 16179 6765
rect 6380 6760 16179 6762
rect 6380 6704 9402 6760
rect 9458 6704 16118 6760
rect 16174 6704 16179 6760
rect 6380 6702 16179 6704
rect 6380 6700 6386 6702
rect 9397 6699 9463 6702
rect 16113 6699 16179 6702
rect 16297 6762 16363 6765
rect 18689 6762 18755 6765
rect 16297 6760 18755 6762
rect 16297 6704 16302 6760
rect 16358 6704 18694 6760
rect 18750 6704 18755 6760
rect 16297 6702 18755 6704
rect 16297 6699 16363 6702
rect 18689 6699 18755 6702
rect 19333 6762 19399 6765
rect 30373 6762 30439 6765
rect 19333 6760 30439 6762
rect 19333 6704 19338 6760
rect 19394 6704 30378 6760
rect 30434 6704 30439 6760
rect 19333 6702 30439 6704
rect 19333 6699 19399 6702
rect 30373 6699 30439 6702
rect 3601 6626 3667 6629
rect 14273 6626 14339 6629
rect 17585 6626 17651 6629
rect 18505 6626 18571 6629
rect 3601 6624 14339 6626
rect 3601 6568 3606 6624
rect 3662 6568 14278 6624
rect 14334 6568 14339 6624
rect 3601 6566 14339 6568
rect 3601 6563 3667 6566
rect 14273 6563 14339 6566
rect 14414 6566 15394 6626
rect 7189 6492 7255 6493
rect 7189 6490 7236 6492
rect 7144 6488 7236 6490
rect 7144 6432 7194 6488
rect 7144 6430 7236 6432
rect 7189 6428 7236 6430
rect 7300 6428 7306 6492
rect 12893 6490 12959 6493
rect 14414 6490 14474 6566
rect 12893 6488 14474 6490
rect 12893 6432 12898 6488
rect 12954 6432 14474 6488
rect 12893 6430 14474 6432
rect 14917 6490 14983 6493
rect 15142 6490 15148 6492
rect 14917 6488 15148 6490
rect 14917 6432 14922 6488
rect 14978 6432 15148 6488
rect 14917 6430 15148 6432
rect 7189 6427 7255 6428
rect 12893 6427 12959 6430
rect 14917 6427 14983 6430
rect 15142 6428 15148 6430
rect 15212 6428 15218 6492
rect 15334 6490 15394 6566
rect 17585 6624 18571 6626
rect 17585 6568 17590 6624
rect 17646 6568 18510 6624
rect 18566 6568 18571 6624
rect 17585 6566 18571 6568
rect 17585 6563 17651 6566
rect 18505 6563 18571 6566
rect 19977 6626 20043 6629
rect 23933 6626 23999 6629
rect 19977 6624 23999 6626
rect 19977 6568 19982 6624
rect 20038 6568 23938 6624
rect 23994 6568 23999 6624
rect 19977 6566 23999 6568
rect 19977 6563 20043 6566
rect 23933 6563 23999 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 19374 6490 19380 6492
rect 15334 6430 19380 6490
rect 19374 6428 19380 6430
rect 19444 6428 19450 6492
rect 1945 6354 2011 6357
rect 24669 6354 24735 6357
rect 1945 6352 24735 6354
rect 1945 6296 1950 6352
rect 2006 6296 24674 6352
rect 24730 6296 24735 6352
rect 1945 6294 24735 6296
rect 1945 6291 2011 6294
rect 24669 6291 24735 6294
rect 4613 6218 4679 6221
rect 8569 6218 8635 6221
rect 4613 6216 8635 6218
rect 4613 6160 4618 6216
rect 4674 6160 8574 6216
rect 8630 6160 8635 6216
rect 4613 6158 8635 6160
rect 4613 6155 4679 6158
rect 8569 6155 8635 6158
rect 13537 6218 13603 6221
rect 13670 6218 13676 6220
rect 13537 6216 13676 6218
rect 13537 6160 13542 6216
rect 13598 6160 13676 6216
rect 13537 6158 13676 6160
rect 13537 6155 13603 6158
rect 13670 6156 13676 6158
rect 13740 6156 13746 6220
rect 16113 6218 16179 6221
rect 23565 6218 23631 6221
rect 16113 6216 23631 6218
rect 16113 6160 16118 6216
rect 16174 6160 23570 6216
rect 23626 6160 23631 6216
rect 16113 6158 23631 6160
rect 16113 6155 16179 6158
rect 23565 6155 23631 6158
rect 38285 6218 38351 6221
rect 39200 6218 39800 6248
rect 38285 6216 39800 6218
rect 38285 6160 38290 6216
rect 38346 6160 39800 6216
rect 38285 6158 39800 6160
rect 38285 6155 38351 6158
rect 39200 6128 39800 6158
rect 7189 6082 7255 6085
rect 12617 6082 12683 6085
rect 21817 6082 21883 6085
rect 7189 6080 12683 6082
rect 7189 6024 7194 6080
rect 7250 6024 12622 6080
rect 12678 6024 12683 6080
rect 7189 6022 12683 6024
rect 7189 6019 7255 6022
rect 12617 6019 12683 6022
rect 13862 6080 21883 6082
rect 13862 6024 21822 6080
rect 21878 6024 21883 6080
rect 13862 6022 21883 6024
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 13261 5946 13327 5949
rect 13862 5946 13922 6022
rect 21817 6019 21883 6022
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 13261 5944 13922 5946
rect 13261 5888 13266 5944
rect 13322 5888 13922 5944
rect 13261 5886 13922 5888
rect 16481 5946 16547 5949
rect 21265 5946 21331 5949
rect 16481 5944 21331 5946
rect 16481 5888 16486 5944
rect 16542 5888 21270 5944
rect 21326 5888 21331 5944
rect 16481 5886 21331 5888
rect 13261 5883 13327 5886
rect 16481 5883 16547 5886
rect 21265 5883 21331 5886
rect 10501 5810 10567 5813
rect 13537 5810 13603 5813
rect 10501 5808 13603 5810
rect 10501 5752 10506 5808
rect 10562 5752 13542 5808
rect 13598 5752 13603 5808
rect 10501 5750 13603 5752
rect 10501 5747 10567 5750
rect 13537 5747 13603 5750
rect 16573 5810 16639 5813
rect 21173 5810 21239 5813
rect 16573 5808 21239 5810
rect 16573 5752 16578 5808
rect 16634 5752 21178 5808
rect 21234 5752 21239 5808
rect 16573 5750 21239 5752
rect 16573 5747 16639 5750
rect 21173 5747 21239 5750
rect 21357 5810 21423 5813
rect 28165 5810 28231 5813
rect 21357 5808 28231 5810
rect 21357 5752 21362 5808
rect 21418 5752 28170 5808
rect 28226 5752 28231 5808
rect 21357 5750 28231 5752
rect 21357 5747 21423 5750
rect 28165 5747 28231 5750
rect 10869 5674 10935 5677
rect 12617 5674 12683 5677
rect 13261 5674 13327 5677
rect 10869 5672 12450 5674
rect 10869 5616 10874 5672
rect 10930 5616 12450 5672
rect 10869 5614 12450 5616
rect 10869 5611 10935 5614
rect 200 5538 800 5568
rect 9949 5538 10015 5541
rect 12249 5538 12315 5541
rect 200 5448 858 5538
rect 9949 5536 12315 5538
rect 9949 5480 9954 5536
rect 10010 5480 12254 5536
rect 12310 5480 12315 5536
rect 9949 5478 12315 5480
rect 12390 5538 12450 5614
rect 12617 5672 13327 5674
rect 12617 5616 12622 5672
rect 12678 5616 13266 5672
rect 13322 5616 13327 5672
rect 12617 5614 13327 5616
rect 12617 5611 12683 5614
rect 13261 5611 13327 5614
rect 15285 5674 15351 5677
rect 18689 5674 18755 5677
rect 15285 5672 18755 5674
rect 15285 5616 15290 5672
rect 15346 5616 18694 5672
rect 18750 5616 18755 5672
rect 15285 5614 18755 5616
rect 15285 5611 15351 5614
rect 18689 5611 18755 5614
rect 19517 5674 19583 5677
rect 21633 5674 21699 5677
rect 19517 5672 21699 5674
rect 19517 5616 19522 5672
rect 19578 5616 21638 5672
rect 21694 5616 21699 5672
rect 19517 5614 21699 5616
rect 19517 5611 19583 5614
rect 21633 5611 21699 5614
rect 21817 5674 21883 5677
rect 23289 5674 23355 5677
rect 21817 5672 23355 5674
rect 21817 5616 21822 5672
rect 21878 5616 23294 5672
rect 23350 5616 23355 5672
rect 21817 5614 23355 5616
rect 21817 5611 21883 5614
rect 23289 5611 23355 5614
rect 13905 5538 13971 5541
rect 12390 5536 13971 5538
rect 12390 5480 13910 5536
rect 13966 5480 13971 5536
rect 12390 5478 13971 5480
rect 9949 5475 10015 5478
rect 12249 5475 12315 5478
rect 13905 5475 13971 5478
rect 16021 5538 16087 5541
rect 19149 5538 19215 5541
rect 16021 5536 19215 5538
rect 16021 5480 16026 5536
rect 16082 5480 19154 5536
rect 19210 5480 19215 5536
rect 16021 5478 19215 5480
rect 16021 5475 16087 5478
rect 19149 5475 19215 5478
rect 20437 5538 20503 5541
rect 22093 5538 22159 5541
rect 20437 5536 22159 5538
rect 20437 5480 20442 5536
rect 20498 5480 22098 5536
rect 22154 5480 22159 5536
rect 20437 5478 22159 5480
rect 20437 5475 20503 5478
rect 22093 5475 22159 5478
rect 798 5266 858 5448
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 9857 5402 9923 5405
rect 15377 5402 15443 5405
rect 9857 5400 15443 5402
rect 9857 5344 9862 5400
rect 9918 5344 15382 5400
rect 15438 5344 15443 5400
rect 9857 5342 15443 5344
rect 9857 5339 9923 5342
rect 15377 5339 15443 5342
rect 17401 5402 17467 5405
rect 19241 5402 19307 5405
rect 17401 5400 19307 5402
rect 17401 5344 17406 5400
rect 17462 5344 19246 5400
rect 19302 5344 19307 5400
rect 17401 5342 19307 5344
rect 17401 5339 17467 5342
rect 19241 5339 19307 5342
rect 20161 5402 20227 5405
rect 20897 5402 20963 5405
rect 20161 5400 20963 5402
rect 20161 5344 20166 5400
rect 20222 5344 20902 5400
rect 20958 5344 20963 5400
rect 20161 5342 20963 5344
rect 20161 5339 20227 5342
rect 20897 5339 20963 5342
rect 21265 5402 21331 5405
rect 21725 5402 21791 5405
rect 21265 5400 21791 5402
rect 21265 5344 21270 5400
rect 21326 5344 21730 5400
rect 21786 5344 21791 5400
rect 21265 5342 21791 5344
rect 21265 5339 21331 5342
rect 21725 5339 21791 5342
rect 614 5206 858 5266
rect 4429 5266 4495 5269
rect 6913 5266 6979 5269
rect 4429 5264 6979 5266
rect 4429 5208 4434 5264
rect 4490 5208 6918 5264
rect 6974 5208 6979 5264
rect 4429 5206 6979 5208
rect 614 4858 674 5206
rect 4429 5203 4495 5206
rect 6913 5203 6979 5206
rect 12065 5266 12131 5269
rect 12341 5266 12407 5269
rect 17585 5266 17651 5269
rect 25865 5266 25931 5269
rect 12065 5264 17418 5266
rect 12065 5208 12070 5264
rect 12126 5208 12346 5264
rect 12402 5208 17418 5264
rect 12065 5206 17418 5208
rect 12065 5203 12131 5206
rect 12341 5203 12407 5206
rect 2681 5130 2747 5133
rect 5717 5130 5783 5133
rect 2681 5128 5783 5130
rect 2681 5072 2686 5128
rect 2742 5072 5722 5128
rect 5778 5072 5783 5128
rect 2681 5070 5783 5072
rect 2681 5067 2747 5070
rect 5717 5067 5783 5070
rect 11973 5130 12039 5133
rect 17358 5130 17418 5206
rect 17585 5264 25931 5266
rect 17585 5208 17590 5264
rect 17646 5208 25870 5264
rect 25926 5208 25931 5264
rect 17585 5206 25931 5208
rect 17585 5203 17651 5206
rect 25865 5203 25931 5206
rect 21081 5130 21147 5133
rect 22737 5130 22803 5133
rect 11973 5128 14290 5130
rect 11973 5072 11978 5128
rect 12034 5072 14290 5128
rect 11973 5070 14290 5072
rect 17358 5128 22803 5130
rect 17358 5072 21086 5128
rect 21142 5072 22742 5128
rect 22798 5072 22803 5128
rect 17358 5070 22803 5072
rect 11973 5067 12039 5070
rect 7741 4994 7807 4997
rect 14089 4994 14155 4997
rect 7741 4992 14155 4994
rect 7741 4936 7746 4992
rect 7802 4936 14094 4992
rect 14150 4936 14155 4992
rect 7741 4934 14155 4936
rect 14230 4994 14290 5070
rect 21081 5067 21147 5070
rect 22737 5067 22803 5070
rect 17401 4994 17467 4997
rect 14230 4992 17467 4994
rect 14230 4936 17406 4992
rect 17462 4936 17467 4992
rect 14230 4934 17467 4936
rect 7741 4931 7807 4934
rect 14089 4931 14155 4934
rect 17401 4931 17467 4934
rect 17769 4994 17835 4997
rect 19149 4994 19215 4997
rect 17769 4992 19215 4994
rect 17769 4936 17774 4992
rect 17830 4936 19154 4992
rect 19210 4936 19215 4992
rect 17769 4934 19215 4936
rect 17769 4931 17835 4934
rect 19149 4931 19215 4934
rect 19425 4994 19491 4997
rect 22001 4994 22067 4997
rect 19425 4992 22067 4994
rect 19425 4936 19430 4992
rect 19486 4936 22006 4992
rect 22062 4936 22067 4992
rect 19425 4934 22067 4936
rect 19425 4931 19491 4934
rect 22001 4931 22067 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 13486 4858 13492 4860
rect 614 4798 2790 4858
rect 2730 4722 2790 4798
rect 4662 4798 13492 4858
rect 4662 4722 4722 4798
rect 13486 4796 13492 4798
rect 13556 4796 13562 4860
rect 13997 4858 14063 4861
rect 17309 4858 17375 4861
rect 13997 4856 17375 4858
rect 13997 4800 14002 4856
rect 14058 4800 17314 4856
rect 17370 4800 17375 4856
rect 13997 4798 17375 4800
rect 13997 4795 14063 4798
rect 17309 4795 17375 4798
rect 17677 4858 17743 4861
rect 23381 4858 23447 4861
rect 17677 4856 23447 4858
rect 17677 4800 17682 4856
rect 17738 4800 23386 4856
rect 23442 4800 23447 4856
rect 17677 4798 23447 4800
rect 17677 4795 17743 4798
rect 23381 4795 23447 4798
rect 38193 4858 38259 4861
rect 39200 4858 39800 4888
rect 38193 4856 39800 4858
rect 38193 4800 38198 4856
rect 38254 4800 39800 4856
rect 38193 4798 39800 4800
rect 38193 4795 38259 4798
rect 39200 4768 39800 4798
rect 2730 4662 4722 4722
rect 10041 4722 10107 4725
rect 22001 4722 22067 4725
rect 10041 4720 22067 4722
rect 10041 4664 10046 4720
rect 10102 4664 22006 4720
rect 22062 4664 22067 4720
rect 10041 4662 22067 4664
rect 10041 4659 10107 4662
rect 22001 4659 22067 4662
rect 5717 4586 5783 4589
rect 6310 4586 6316 4588
rect 5717 4584 6316 4586
rect 5717 4528 5722 4584
rect 5778 4528 6316 4584
rect 5717 4526 6316 4528
rect 5717 4523 5783 4526
rect 6310 4524 6316 4526
rect 6380 4524 6386 4588
rect 12157 4586 12223 4589
rect 12525 4586 12591 4589
rect 12157 4584 12591 4586
rect 12157 4528 12162 4584
rect 12218 4528 12530 4584
rect 12586 4528 12591 4584
rect 12157 4526 12591 4528
rect 12157 4523 12223 4526
rect 12525 4523 12591 4526
rect 14273 4586 14339 4589
rect 20437 4586 20503 4589
rect 23657 4586 23723 4589
rect 14273 4584 20132 4586
rect 14273 4528 14278 4584
rect 14334 4528 20132 4584
rect 14273 4526 20132 4528
rect 14273 4523 14339 4526
rect 12065 4450 12131 4453
rect 12341 4450 12407 4453
rect 12065 4448 12407 4450
rect 12065 4392 12070 4448
rect 12126 4392 12346 4448
rect 12402 4392 12407 4448
rect 12065 4390 12407 4392
rect 12065 4387 12131 4390
rect 12341 4387 12407 4390
rect 13537 4450 13603 4453
rect 16021 4450 16087 4453
rect 13537 4448 16087 4450
rect 13537 4392 13542 4448
rect 13598 4392 16026 4448
rect 16082 4392 16087 4448
rect 13537 4390 16087 4392
rect 20072 4450 20132 4526
rect 20437 4584 23723 4586
rect 20437 4528 20442 4584
rect 20498 4528 23662 4584
rect 23718 4528 23723 4584
rect 20437 4526 23723 4528
rect 20437 4523 20503 4526
rect 23657 4523 23723 4526
rect 25497 4450 25563 4453
rect 20072 4448 25563 4450
rect 20072 4392 25502 4448
rect 25558 4392 25563 4448
rect 20072 4390 25563 4392
rect 13537 4387 13603 4390
rect 16021 4387 16087 4390
rect 25497 4387 25563 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4705 4314 4771 4317
rect 5073 4314 5139 4317
rect 4705 4312 5139 4314
rect 4705 4256 4710 4312
rect 4766 4256 5078 4312
rect 5134 4256 5139 4312
rect 4705 4254 5139 4256
rect 4705 4251 4771 4254
rect 5073 4251 5139 4254
rect 11145 4314 11211 4317
rect 18321 4314 18387 4317
rect 20161 4316 20227 4317
rect 11145 4312 18387 4314
rect 11145 4256 11150 4312
rect 11206 4256 18326 4312
rect 18382 4256 18387 4312
rect 11145 4254 18387 4256
rect 11145 4251 11211 4254
rect 18321 4251 18387 4254
rect 20110 4252 20116 4316
rect 20180 4314 20227 4316
rect 20897 4314 20963 4317
rect 22737 4314 22803 4317
rect 20180 4312 20272 4314
rect 20222 4256 20272 4312
rect 20180 4254 20272 4256
rect 20897 4312 22803 4314
rect 20897 4256 20902 4312
rect 20958 4256 22742 4312
rect 22798 4256 22803 4312
rect 20897 4254 22803 4256
rect 20180 4252 20227 4254
rect 20161 4251 20227 4252
rect 20897 4251 20963 4254
rect 22737 4251 22803 4254
rect 200 4178 800 4208
rect 1761 4178 1827 4181
rect 200 4176 1827 4178
rect 200 4120 1766 4176
rect 1822 4120 1827 4176
rect 200 4118 1827 4120
rect 200 4088 800 4118
rect 1761 4115 1827 4118
rect 7373 4178 7439 4181
rect 15377 4178 15443 4181
rect 7373 4176 15443 4178
rect 7373 4120 7378 4176
rect 7434 4120 15382 4176
rect 15438 4120 15443 4176
rect 7373 4118 15443 4120
rect 7373 4115 7439 4118
rect 15377 4115 15443 4118
rect 15745 4178 15811 4181
rect 17677 4178 17743 4181
rect 15745 4176 17743 4178
rect 15745 4120 15750 4176
rect 15806 4120 17682 4176
rect 17738 4120 17743 4176
rect 15745 4118 17743 4120
rect 15745 4115 15811 4118
rect 17677 4115 17743 4118
rect 19333 4178 19399 4181
rect 20713 4178 20779 4181
rect 19333 4176 20779 4178
rect 19333 4120 19338 4176
rect 19394 4120 20718 4176
rect 20774 4120 20779 4176
rect 19333 4118 20779 4120
rect 19333 4115 19399 4118
rect 20713 4115 20779 4118
rect 38285 4178 38351 4181
rect 39200 4178 39800 4208
rect 38285 4176 39800 4178
rect 38285 4120 38290 4176
rect 38346 4120 39800 4176
rect 38285 4118 39800 4120
rect 38285 4115 38351 4118
rect 39200 4088 39800 4118
rect 4521 4042 4587 4045
rect 5073 4042 5139 4045
rect 4521 4040 5139 4042
rect 4521 3984 4526 4040
rect 4582 3984 5078 4040
rect 5134 3984 5139 4040
rect 4521 3982 5139 3984
rect 4521 3979 4587 3982
rect 5073 3979 5139 3982
rect 6729 4042 6795 4045
rect 13445 4042 13511 4045
rect 6729 4040 13511 4042
rect 6729 3984 6734 4040
rect 6790 3984 13450 4040
rect 13506 3984 13511 4040
rect 6729 3982 13511 3984
rect 6729 3979 6795 3982
rect 13445 3979 13511 3982
rect 13905 4042 13971 4045
rect 20529 4042 20595 4045
rect 13905 4040 20595 4042
rect 13905 3984 13910 4040
rect 13966 3984 20534 4040
rect 20590 3984 20595 4040
rect 13905 3982 20595 3984
rect 13905 3979 13971 3982
rect 20529 3979 20595 3982
rect 9397 3906 9463 3909
rect 11513 3906 11579 3909
rect 12157 3906 12223 3909
rect 15009 3906 15075 3909
rect 9397 3904 12223 3906
rect 9397 3848 9402 3904
rect 9458 3848 11518 3904
rect 11574 3848 12162 3904
rect 12218 3848 12223 3904
rect 9397 3846 12223 3848
rect 9397 3843 9463 3846
rect 11513 3843 11579 3846
rect 12157 3843 12223 3846
rect 12390 3904 15075 3906
rect 12390 3848 15014 3904
rect 15070 3848 15075 3904
rect 12390 3846 15075 3848
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12390 3770 12450 3846
rect 15009 3843 15075 3846
rect 17677 3906 17743 3909
rect 22829 3906 22895 3909
rect 17677 3904 22895 3906
rect 17677 3848 17682 3904
rect 17738 3848 22834 3904
rect 22890 3848 22895 3904
rect 17677 3846 22895 3848
rect 17677 3843 17743 3846
rect 22829 3843 22895 3846
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 6318 3710 12450 3770
rect 14181 3770 14247 3773
rect 23289 3770 23355 3773
rect 14181 3768 23355 3770
rect 14181 3712 14186 3768
rect 14242 3712 23294 3768
rect 23350 3712 23355 3768
rect 14181 3710 23355 3712
rect 4337 3634 4403 3637
rect 6318 3634 6378 3710
rect 14181 3707 14247 3710
rect 23289 3707 23355 3710
rect 4337 3632 6378 3634
rect 4337 3576 4342 3632
rect 4398 3576 6378 3632
rect 4337 3574 6378 3576
rect 4337 3571 4403 3574
rect 6678 3572 6684 3636
rect 6748 3634 6754 3636
rect 6821 3634 6887 3637
rect 6748 3632 6887 3634
rect 6748 3576 6826 3632
rect 6882 3576 6887 3632
rect 6748 3574 6887 3576
rect 6748 3572 6754 3574
rect 6821 3571 6887 3574
rect 14365 3634 14431 3637
rect 15837 3634 15903 3637
rect 14365 3632 15903 3634
rect 14365 3576 14370 3632
rect 14426 3576 15842 3632
rect 15898 3576 15903 3632
rect 14365 3574 15903 3576
rect 14365 3571 14431 3574
rect 15837 3571 15903 3574
rect 16481 3634 16547 3637
rect 21817 3634 21883 3637
rect 16481 3632 21883 3634
rect 16481 3576 16486 3632
rect 16542 3576 21822 3632
rect 21878 3576 21883 3632
rect 16481 3574 21883 3576
rect 16481 3571 16547 3574
rect 21817 3571 21883 3574
rect 22093 3634 22159 3637
rect 27981 3634 28047 3637
rect 22093 3632 28047 3634
rect 22093 3576 22098 3632
rect 22154 3576 27986 3632
rect 28042 3576 28047 3632
rect 22093 3574 28047 3576
rect 22093 3571 22159 3574
rect 27981 3571 28047 3574
rect 200 3498 800 3528
rect 4061 3498 4127 3501
rect 200 3496 4127 3498
rect 200 3440 4066 3496
rect 4122 3440 4127 3496
rect 200 3438 4127 3440
rect 200 3408 800 3438
rect 4061 3435 4127 3438
rect 4337 3498 4403 3501
rect 6545 3498 6611 3501
rect 4337 3496 6611 3498
rect 4337 3440 4342 3496
rect 4398 3440 6550 3496
rect 6606 3440 6611 3496
rect 4337 3438 6611 3440
rect 4337 3435 4403 3438
rect 6545 3435 6611 3438
rect 10225 3498 10291 3501
rect 11973 3498 12039 3501
rect 27797 3498 27863 3501
rect 10225 3496 12039 3498
rect 10225 3440 10230 3496
rect 10286 3440 11978 3496
rect 12034 3440 12039 3496
rect 10225 3438 12039 3440
rect 10225 3435 10291 3438
rect 11973 3435 12039 3438
rect 12390 3496 27863 3498
rect 12390 3440 27802 3496
rect 27858 3440 27863 3496
rect 12390 3438 27863 3440
rect 1577 3362 1643 3365
rect 12390 3362 12450 3438
rect 27797 3435 27863 3438
rect 1577 3360 12450 3362
rect 1577 3304 1582 3360
rect 1638 3304 12450 3360
rect 1577 3302 12450 3304
rect 15193 3362 15259 3365
rect 16389 3362 16455 3365
rect 15193 3360 16455 3362
rect 15193 3304 15198 3360
rect 15254 3304 16394 3360
rect 16450 3304 16455 3360
rect 15193 3302 16455 3304
rect 1577 3299 1643 3302
rect 15193 3299 15259 3302
rect 16389 3299 16455 3302
rect 20069 3362 20135 3365
rect 20529 3362 20595 3365
rect 20069 3360 20595 3362
rect 20069 3304 20074 3360
rect 20130 3304 20534 3360
rect 20590 3304 20595 3360
rect 20069 3302 20595 3304
rect 20069 3299 20135 3302
rect 20529 3299 20595 3302
rect 20713 3362 20779 3365
rect 26601 3362 26667 3365
rect 20713 3360 26667 3362
rect 20713 3304 20718 3360
rect 20774 3304 26606 3360
rect 26662 3304 26667 3360
rect 20713 3302 26667 3304
rect 20713 3299 20779 3302
rect 26601 3299 26667 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 5809 3226 5875 3229
rect 7833 3226 7899 3229
rect 5809 3224 7899 3226
rect 5809 3168 5814 3224
rect 5870 3168 7838 3224
rect 7894 3168 7899 3224
rect 5809 3166 7899 3168
rect 5809 3163 5875 3166
rect 7833 3163 7899 3166
rect 8017 3226 8083 3229
rect 16021 3226 16087 3229
rect 8017 3224 16087 3226
rect 8017 3168 8022 3224
rect 8078 3168 16026 3224
rect 16082 3168 16087 3224
rect 8017 3166 16087 3168
rect 8017 3163 8083 3166
rect 16021 3163 16087 3166
rect 20161 3226 20227 3229
rect 22645 3226 22711 3229
rect 20161 3224 22711 3226
rect 20161 3168 20166 3224
rect 20222 3168 22650 3224
rect 22706 3168 22711 3224
rect 20161 3166 22711 3168
rect 20161 3163 20227 3166
rect 22645 3163 22711 3166
rect 5073 3090 5139 3093
rect 19609 3090 19675 3093
rect 5073 3088 19675 3090
rect 5073 3032 5078 3088
rect 5134 3032 19614 3088
rect 19670 3032 19675 3088
rect 5073 3030 19675 3032
rect 5073 3027 5139 3030
rect 19609 3027 19675 3030
rect 19977 3090 20043 3093
rect 22461 3090 22527 3093
rect 19977 3088 22527 3090
rect 19977 3032 19982 3088
rect 20038 3032 22466 3088
rect 22522 3032 22527 3088
rect 19977 3030 22527 3032
rect 19977 3027 20043 3030
rect 22461 3027 22527 3030
rect 5165 2954 5231 2957
rect 7373 2954 7439 2957
rect 5165 2952 7439 2954
rect 5165 2896 5170 2952
rect 5226 2896 7378 2952
rect 7434 2896 7439 2952
rect 5165 2894 7439 2896
rect 5165 2891 5231 2894
rect 7373 2891 7439 2894
rect 14457 2954 14523 2957
rect 20161 2954 20227 2957
rect 20345 2956 20411 2957
rect 14457 2952 20227 2954
rect 14457 2896 14462 2952
rect 14518 2896 20166 2952
rect 20222 2896 20227 2952
rect 14457 2894 20227 2896
rect 14457 2891 14523 2894
rect 20161 2891 20227 2894
rect 20294 2892 20300 2956
rect 20364 2954 20411 2956
rect 21909 2954 21975 2957
rect 20364 2952 20456 2954
rect 20406 2896 20456 2952
rect 20364 2894 20456 2896
rect 20670 2952 21975 2954
rect 20670 2896 21914 2952
rect 21970 2896 21975 2952
rect 20670 2894 21975 2896
rect 20364 2892 20411 2894
rect 20345 2891 20411 2892
rect 9673 2818 9739 2821
rect 10593 2818 10659 2821
rect 14917 2818 14983 2821
rect 9673 2816 14983 2818
rect 9673 2760 9678 2816
rect 9734 2760 10598 2816
rect 10654 2760 14922 2816
rect 14978 2760 14983 2816
rect 9673 2758 14983 2760
rect 9673 2755 9739 2758
rect 10593 2755 10659 2758
rect 14917 2755 14983 2758
rect 19057 2818 19123 2821
rect 20670 2818 20730 2894
rect 21909 2891 21975 2894
rect 19057 2816 20730 2818
rect 19057 2760 19062 2816
rect 19118 2760 20730 2816
rect 19057 2758 20730 2760
rect 21633 2818 21699 2821
rect 22553 2818 22619 2821
rect 21633 2816 22619 2818
rect 21633 2760 21638 2816
rect 21694 2760 22558 2816
rect 22614 2760 22619 2816
rect 21633 2758 22619 2760
rect 19057 2755 19123 2758
rect 21633 2755 21699 2758
rect 22553 2755 22619 2758
rect 38193 2818 38259 2821
rect 39200 2818 39800 2848
rect 38193 2816 39800 2818
rect 38193 2760 38198 2816
rect 38254 2760 39800 2816
rect 38193 2758 39800 2760
rect 38193 2755 38259 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 3141 2684 3207 2685
rect 15377 2684 15443 2685
rect 3141 2680 3188 2684
rect 3252 2682 3258 2684
rect 3141 2624 3146 2680
rect 3141 2620 3188 2624
rect 3252 2622 3298 2682
rect 3252 2620 3258 2622
rect 15326 2620 15332 2684
rect 15396 2682 15443 2684
rect 17217 2682 17283 2685
rect 22737 2682 22803 2685
rect 15396 2680 15488 2682
rect 15438 2624 15488 2680
rect 15396 2622 15488 2624
rect 17217 2680 22803 2682
rect 17217 2624 17222 2680
rect 17278 2624 22742 2680
rect 22798 2624 22803 2680
rect 17217 2622 22803 2624
rect 15396 2620 15443 2622
rect 3141 2619 3207 2620
rect 15377 2619 15443 2620
rect 17217 2619 17283 2622
rect 22737 2619 22803 2622
rect 3877 2546 3943 2549
rect 23381 2546 23447 2549
rect 3877 2544 23447 2546
rect 3877 2488 3882 2544
rect 3938 2488 23386 2544
rect 23442 2488 23447 2544
rect 3877 2486 23447 2488
rect 3877 2483 3943 2486
rect 23381 2483 23447 2486
rect 4061 2410 4127 2413
rect 23381 2410 23447 2413
rect 4061 2408 23447 2410
rect 4061 2352 4066 2408
rect 4122 2352 23386 2408
rect 23442 2352 23447 2408
rect 4061 2350 23447 2352
rect 4061 2347 4127 2350
rect 23381 2347 23447 2350
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 1761 2138 1827 2141
rect 200 2136 1827 2138
rect 200 2080 1766 2136
rect 1822 2080 1827 2136
rect 200 2078 1827 2080
rect 200 2048 800 2078
rect 1761 2075 1827 2078
rect 6545 2002 6611 2005
rect 27153 2002 27219 2005
rect 6545 2000 27219 2002
rect 6545 1944 6550 2000
rect 6606 1944 27158 2000
rect 27214 1944 27219 2000
rect 6545 1942 27219 1944
rect 6545 1939 6611 1942
rect 27153 1939 27219 1942
rect 5257 1866 5323 1869
rect 22093 1866 22159 1869
rect 5257 1864 22159 1866
rect 5257 1808 5262 1864
rect 5318 1808 22098 1864
rect 22154 1808 22159 1864
rect 5257 1806 22159 1808
rect 5257 1803 5323 1806
rect 22093 1803 22159 1806
rect 14089 1730 14155 1733
rect 23933 1730 23999 1733
rect 14089 1728 23999 1730
rect 14089 1672 14094 1728
rect 14150 1672 23938 1728
rect 23994 1672 23999 1728
rect 14089 1670 23999 1672
rect 14089 1667 14155 1670
rect 23933 1667 23999 1670
rect 3693 1594 3759 1597
rect 24025 1594 24091 1597
rect 3693 1592 24091 1594
rect 3693 1536 3698 1592
rect 3754 1536 24030 1592
rect 24086 1536 24091 1592
rect 3693 1534 24091 1536
rect 3693 1531 3759 1534
rect 24025 1531 24091 1534
rect 37181 1458 37247 1461
rect 39200 1458 39800 1488
rect 37181 1456 39800 1458
rect 37181 1400 37186 1456
rect 37242 1400 39800 1456
rect 37181 1398 39800 1400
rect 37181 1395 37247 1398
rect 39200 1368 39800 1398
rect 200 778 800 808
rect 1393 778 1459 781
rect 200 776 1459 778
rect 200 720 1398 776
rect 1454 720 1459 776
rect 200 718 1459 720
rect 200 688 800 718
rect 1393 715 1459 718
rect 37457 778 37523 781
rect 39200 778 39800 808
rect 37457 776 39800 778
rect 37457 720 37462 776
rect 37518 720 39800 776
rect 37457 718 39800 720
rect 37457 715 37523 718
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 2452 35940 2516 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 6132 30364 6196 30428
rect 18092 30228 18156 30292
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 1716 26828 1780 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 2636 26556 2700 26620
rect 1900 26284 1964 26348
rect 3372 26284 3436 26348
rect 6500 26344 6564 26348
rect 6500 26288 6514 26344
rect 6514 26288 6564 26344
rect 6500 26284 6564 26288
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 3740 25604 3804 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 3924 24984 3988 24988
rect 3924 24928 3974 24984
rect 3974 24928 3988 24984
rect 3924 24924 3988 24928
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4660 23972 4724 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 10732 23836 10796 23900
rect 5580 23700 5644 23764
rect 7236 23564 7300 23628
rect 11100 23428 11164 23492
rect 12572 23428 12636 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 15516 22884 15580 22948
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 5948 22808 6012 22812
rect 5948 22752 5998 22808
rect 5998 22752 6012 22808
rect 5948 22748 6012 22752
rect 2820 22612 2884 22676
rect 15516 22612 15580 22676
rect 5764 22536 5828 22540
rect 5764 22480 5778 22536
rect 5778 22480 5828 22536
rect 5764 22476 5828 22480
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 6316 22128 6380 22132
rect 6316 22072 6330 22128
rect 6330 22072 6380 22128
rect 6316 22068 6380 22072
rect 5580 21932 5644 21996
rect 9628 22068 9692 22132
rect 10732 21992 10796 21996
rect 10732 21936 10782 21992
rect 10782 21936 10796 21992
rect 10732 21932 10796 21936
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4660 21524 4724 21588
rect 5948 21252 6012 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 6316 20980 6380 21044
rect 14228 20844 14292 20908
rect 17724 20708 17788 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 2820 20572 2884 20636
rect 3188 20436 3252 20500
rect 12572 20436 12636 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 6132 19816 6196 19820
rect 6132 19760 6182 19816
rect 6182 19760 6196 19816
rect 6132 19756 6196 19760
rect 12940 19756 13004 19820
rect 11100 19620 11164 19684
rect 11652 19620 11716 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 1900 19484 1964 19548
rect 3740 19544 3804 19548
rect 3740 19488 3754 19544
rect 3754 19488 3804 19544
rect 3740 19484 3804 19488
rect 3924 19348 3988 19412
rect 5028 19348 5092 19412
rect 7052 19408 7116 19412
rect 7052 19352 7066 19408
rect 7066 19352 7116 19408
rect 7052 19348 7116 19352
rect 9628 19212 9692 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 12572 18804 12636 18868
rect 6684 18532 6748 18596
rect 14044 18532 14108 18596
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 7236 18260 7300 18324
rect 5764 18048 5828 18052
rect 5764 17992 5778 18048
rect 5778 17992 5828 18048
rect 5764 17988 5828 17992
rect 17356 17988 17420 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 3372 17912 3436 17916
rect 3372 17856 3386 17912
rect 3386 17856 3436 17912
rect 3372 17852 3436 17856
rect 16252 17444 16316 17508
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 1716 17308 1780 17372
rect 20116 17232 20180 17236
rect 20116 17176 20166 17232
rect 20166 17176 20180 17232
rect 20116 17172 20180 17176
rect 3924 16900 3988 16964
rect 9444 16960 9508 16964
rect 9444 16904 9458 16960
rect 9458 16904 9508 16960
rect 9444 16900 9508 16904
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 10916 16688 10980 16692
rect 10916 16632 10966 16688
rect 10966 16632 10980 16688
rect 10916 16628 10980 16632
rect 7236 16552 7300 16556
rect 7236 16496 7250 16552
rect 7250 16496 7300 16552
rect 7236 16492 7300 16496
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 6500 16220 6564 16284
rect 8156 16220 8220 16284
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 12572 15540 12636 15604
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 15516 15192 15580 15196
rect 15516 15136 15530 15192
rect 15530 15136 15580 15192
rect 15516 15132 15580 15136
rect 10732 14860 10796 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 16252 14588 16316 14652
rect 9444 14376 9508 14380
rect 9444 14320 9494 14376
rect 9494 14320 9508 14376
rect 9444 14316 9508 14320
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 14044 13772 14108 13836
rect 14228 13696 14292 13700
rect 14228 13640 14278 13696
rect 14278 13640 14292 13696
rect 14228 13636 14292 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 18092 13500 18156 13564
rect 10916 13092 10980 13156
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 8156 12684 8220 12748
rect 20116 12684 20180 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 1900 11928 1964 11932
rect 1900 11872 1914 11928
rect 1914 11872 1964 11928
rect 1900 11868 1964 11872
rect 3924 11732 3988 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 11652 11188 11716 11252
rect 15148 11188 15212 11252
rect 10732 11052 10796 11116
rect 13676 11052 13740 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 2452 10780 2516 10844
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 17724 10236 17788 10300
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 7052 9692 7116 9756
rect 5028 9420 5092 9484
rect 15332 9420 15396 9484
rect 19380 9420 19444 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 2636 9208 2700 9212
rect 2636 9152 2650 9208
rect 2650 9152 2700 9208
rect 2636 9148 2700 9152
rect 20300 8876 20364 8940
rect 19380 8800 19444 8804
rect 19380 8744 19394 8800
rect 19394 8744 19444 8800
rect 19380 8740 19444 8744
rect 20116 8800 20180 8804
rect 20116 8744 20166 8800
rect 20166 8744 20180 8800
rect 20116 8740 20180 8744
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 12940 8332 13004 8396
rect 19380 8332 19444 8396
rect 8340 8196 8404 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 17724 7576 17788 7580
rect 17724 7520 17738 7576
rect 17738 7520 17788 7576
rect 17724 7516 17788 7520
rect 13492 7108 13556 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 17356 6972 17420 7036
rect 6316 6700 6380 6764
rect 7236 6488 7300 6492
rect 7236 6432 7250 6488
rect 7250 6432 7300 6488
rect 7236 6428 7300 6432
rect 15148 6428 15212 6492
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 19380 6428 19444 6492
rect 13676 6156 13740 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 13492 4796 13556 4860
rect 6316 4524 6380 4588
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 20116 4312 20180 4316
rect 20116 4256 20166 4312
rect 20166 4256 20180 4312
rect 20116 4252 20180 4256
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 6684 3572 6748 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 20300 2952 20364 2956
rect 20300 2896 20350 2952
rect 20350 2896 20364 2952
rect 20300 2892 20364 2896
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 3188 2680 3252 2684
rect 3188 2624 3202 2680
rect 3202 2624 3252 2680
rect 3188 2620 3252 2624
rect 15332 2680 15396 2684
rect 15332 2624 15382 2680
rect 15382 2624 15396 2680
rect 15332 2620 15396 2624
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 2451 36004 2517 36005
rect 2451 35940 2452 36004
rect 2516 35940 2517 36004
rect 2451 35939 2517 35940
rect 1715 26892 1781 26893
rect 1715 26828 1716 26892
rect 1780 26828 1781 26892
rect 1715 26827 1781 26828
rect 1718 17373 1778 26827
rect 1899 26348 1965 26349
rect 1899 26284 1900 26348
rect 1964 26284 1965 26348
rect 1899 26283 1965 26284
rect 1902 19549 1962 26283
rect 1899 19548 1965 19549
rect 1899 19484 1900 19548
rect 1964 19484 1965 19548
rect 1899 19483 1965 19484
rect 1715 17372 1781 17373
rect 1715 17308 1716 17372
rect 1780 17308 1781 17372
rect 1715 17307 1781 17308
rect 1902 11933 1962 19483
rect 1899 11932 1965 11933
rect 1899 11868 1900 11932
rect 1964 11868 1965 11932
rect 1899 11867 1965 11868
rect 2454 10845 2514 35939
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 6131 30428 6197 30429
rect 6131 30364 6132 30428
rect 6196 30364 6197 30428
rect 6131 30363 6197 30364
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 2635 26620 2701 26621
rect 2635 26556 2636 26620
rect 2700 26556 2701 26620
rect 2635 26555 2701 26556
rect 2451 10844 2517 10845
rect 2451 10780 2452 10844
rect 2516 10780 2517 10844
rect 2451 10779 2517 10780
rect 2638 9213 2698 26555
rect 3371 26348 3437 26349
rect 3371 26284 3372 26348
rect 3436 26284 3437 26348
rect 3371 26283 3437 26284
rect 2819 22676 2885 22677
rect 2819 22612 2820 22676
rect 2884 22612 2885 22676
rect 2819 22611 2885 22612
rect 2822 20637 2882 22611
rect 2819 20636 2885 20637
rect 2819 20572 2820 20636
rect 2884 20572 2885 20636
rect 2819 20571 2885 20572
rect 3187 20500 3253 20501
rect 3187 20436 3188 20500
rect 3252 20436 3253 20500
rect 3187 20435 3253 20436
rect 2635 9212 2701 9213
rect 2635 9148 2636 9212
rect 2700 9148 2701 9212
rect 2635 9147 2701 9148
rect 3190 2685 3250 20435
rect 3374 17917 3434 26283
rect 3739 25668 3805 25669
rect 3739 25604 3740 25668
rect 3804 25604 3805 25668
rect 3739 25603 3805 25604
rect 3742 19549 3802 25603
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 3923 24988 3989 24989
rect 3923 24924 3924 24988
rect 3988 24924 3989 24988
rect 3923 24923 3989 24924
rect 3739 19548 3805 19549
rect 3739 19484 3740 19548
rect 3804 19484 3805 19548
rect 3739 19483 3805 19484
rect 3926 19413 3986 24923
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4659 24036 4725 24037
rect 4659 23972 4660 24036
rect 4724 23972 4725 24036
rect 4659 23971 4725 23972
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4662 21589 4722 23971
rect 5579 23764 5645 23765
rect 5579 23700 5580 23764
rect 5644 23700 5645 23764
rect 5579 23699 5645 23700
rect 5582 21997 5642 23699
rect 5947 22812 6013 22813
rect 5947 22748 5948 22812
rect 6012 22748 6013 22812
rect 5947 22747 6013 22748
rect 5763 22540 5829 22541
rect 5763 22476 5764 22540
rect 5828 22476 5829 22540
rect 5763 22475 5829 22476
rect 5579 21996 5645 21997
rect 5579 21932 5580 21996
rect 5644 21932 5645 21996
rect 5579 21931 5645 21932
rect 4659 21588 4725 21589
rect 4659 21524 4660 21588
rect 4724 21524 4725 21588
rect 4659 21523 4725 21524
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3923 19412 3989 19413
rect 3923 19348 3924 19412
rect 3988 19348 3989 19412
rect 3923 19347 3989 19348
rect 4208 19072 4528 20096
rect 5027 19412 5093 19413
rect 5027 19348 5028 19412
rect 5092 19348 5093 19412
rect 5027 19347 5093 19348
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 3371 17916 3437 17917
rect 3371 17852 3372 17916
rect 3436 17852 3437 17916
rect 3371 17851 3437 17852
rect 3923 16964 3989 16965
rect 3923 16900 3924 16964
rect 3988 16900 3989 16964
rect 3923 16899 3989 16900
rect 3926 11797 3986 16899
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 3923 11796 3989 11797
rect 3923 11732 3924 11796
rect 3988 11732 3989 11796
rect 3923 11731 3989 11732
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 5030 9485 5090 19347
rect 5766 18053 5826 22475
rect 5950 21317 6010 22747
rect 5947 21316 6013 21317
rect 5947 21252 5948 21316
rect 6012 21252 6013 21316
rect 5947 21251 6013 21252
rect 6134 19821 6194 30363
rect 18091 30292 18157 30293
rect 18091 30228 18092 30292
rect 18156 30228 18157 30292
rect 18091 30227 18157 30228
rect 6499 26348 6565 26349
rect 6499 26284 6500 26348
rect 6564 26284 6565 26348
rect 6499 26283 6565 26284
rect 6315 22132 6381 22133
rect 6315 22068 6316 22132
rect 6380 22068 6381 22132
rect 6315 22067 6381 22068
rect 6318 21045 6378 22067
rect 6315 21044 6381 21045
rect 6315 20980 6316 21044
rect 6380 20980 6381 21044
rect 6315 20979 6381 20980
rect 6131 19820 6197 19821
rect 6131 19756 6132 19820
rect 6196 19756 6197 19820
rect 6131 19755 6197 19756
rect 5763 18052 5829 18053
rect 5763 17988 5764 18052
rect 5828 17988 5829 18052
rect 5763 17987 5829 17988
rect 5027 9484 5093 9485
rect 5027 9420 5028 9484
rect 5092 9420 5093 9484
rect 5027 9419 5093 9420
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 6318 6765 6378 20979
rect 6502 16285 6562 26283
rect 10731 23900 10797 23901
rect 10731 23836 10732 23900
rect 10796 23836 10797 23900
rect 10731 23835 10797 23836
rect 7235 23628 7301 23629
rect 7235 23564 7236 23628
rect 7300 23564 7301 23628
rect 7235 23563 7301 23564
rect 7051 19412 7117 19413
rect 7051 19348 7052 19412
rect 7116 19348 7117 19412
rect 7051 19347 7117 19348
rect 6683 18596 6749 18597
rect 6683 18532 6684 18596
rect 6748 18532 6749 18596
rect 6683 18531 6749 18532
rect 6499 16284 6565 16285
rect 6499 16220 6500 16284
rect 6564 16220 6565 16284
rect 6499 16219 6565 16220
rect 6315 6764 6381 6765
rect 6315 6700 6316 6764
rect 6380 6700 6381 6764
rect 6315 6699 6381 6700
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 6318 4589 6378 6699
rect 6315 4588 6381 4589
rect 6315 4524 6316 4588
rect 6380 4524 6381 4588
rect 6315 4523 6381 4524
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 6686 3637 6746 18531
rect 7054 9757 7114 19347
rect 7238 18325 7298 23563
rect 9627 22132 9693 22133
rect 9627 22068 9628 22132
rect 9692 22068 9693 22132
rect 9627 22067 9693 22068
rect 9630 19277 9690 22067
rect 10734 21997 10794 23835
rect 11099 23492 11165 23493
rect 11099 23428 11100 23492
rect 11164 23428 11165 23492
rect 11099 23427 11165 23428
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23428 12637 23492
rect 12571 23427 12637 23428
rect 10731 21996 10797 21997
rect 10731 21932 10732 21996
rect 10796 21932 10797 21996
rect 10731 21931 10797 21932
rect 11102 19685 11162 23427
rect 12574 20501 12634 23427
rect 15515 22948 15581 22949
rect 15515 22884 15516 22948
rect 15580 22884 15581 22948
rect 15515 22883 15581 22884
rect 15518 22677 15578 22883
rect 15515 22676 15581 22677
rect 15515 22612 15516 22676
rect 15580 22612 15581 22676
rect 15515 22611 15581 22612
rect 14227 20908 14293 20909
rect 14227 20844 14228 20908
rect 14292 20844 14293 20908
rect 14227 20843 14293 20844
rect 12571 20500 12637 20501
rect 12571 20436 12572 20500
rect 12636 20436 12637 20500
rect 12571 20435 12637 20436
rect 12939 19820 13005 19821
rect 12939 19756 12940 19820
rect 13004 19756 13005 19820
rect 12939 19755 13005 19756
rect 11099 19684 11165 19685
rect 11099 19620 11100 19684
rect 11164 19620 11165 19684
rect 11099 19619 11165 19620
rect 11651 19684 11717 19685
rect 11651 19620 11652 19684
rect 11716 19620 11717 19684
rect 11651 19619 11717 19620
rect 9627 19276 9693 19277
rect 9627 19212 9628 19276
rect 9692 19212 9693 19276
rect 9627 19211 9693 19212
rect 7235 18324 7301 18325
rect 7235 18260 7236 18324
rect 7300 18260 7301 18324
rect 7235 18259 7301 18260
rect 9443 16964 9509 16965
rect 9443 16900 9444 16964
rect 9508 16900 9509 16964
rect 9443 16899 9509 16900
rect 7235 16556 7301 16557
rect 7235 16492 7236 16556
rect 7300 16492 7301 16556
rect 7235 16491 7301 16492
rect 7051 9756 7117 9757
rect 7051 9692 7052 9756
rect 7116 9692 7117 9756
rect 7051 9691 7117 9692
rect 7238 6493 7298 16491
rect 8155 16284 8221 16285
rect 8155 16220 8156 16284
rect 8220 16220 8221 16284
rect 8155 16219 8221 16220
rect 8158 12749 8218 16219
rect 9446 14381 9506 16899
rect 10915 16692 10981 16693
rect 10915 16628 10916 16692
rect 10980 16628 10981 16692
rect 10915 16627 10981 16628
rect 10731 14924 10797 14925
rect 10731 14860 10732 14924
rect 10796 14860 10797 14924
rect 10731 14859 10797 14860
rect 9443 14380 9509 14381
rect 9443 14316 9444 14380
rect 9508 14316 9509 14380
rect 9443 14315 9509 14316
rect 8155 12748 8221 12749
rect 8155 12684 8156 12748
rect 8220 12684 8221 12748
rect 8155 12683 8221 12684
rect 8158 12450 8218 12683
rect 8158 12390 8402 12450
rect 8342 8261 8402 12390
rect 10734 11117 10794 14859
rect 10918 13157 10978 16627
rect 10915 13156 10981 13157
rect 10915 13092 10916 13156
rect 10980 13092 10981 13156
rect 10915 13091 10981 13092
rect 11654 11253 11714 19619
rect 12571 18868 12637 18869
rect 12571 18804 12572 18868
rect 12636 18804 12637 18868
rect 12571 18803 12637 18804
rect 12574 15605 12634 18803
rect 12571 15604 12637 15605
rect 12571 15540 12572 15604
rect 12636 15540 12637 15604
rect 12571 15539 12637 15540
rect 11651 11252 11717 11253
rect 11651 11188 11652 11252
rect 11716 11188 11717 11252
rect 11651 11187 11717 11188
rect 10731 11116 10797 11117
rect 10731 11052 10732 11116
rect 10796 11052 10797 11116
rect 10731 11051 10797 11052
rect 12942 8397 13002 19755
rect 14043 18596 14109 18597
rect 14043 18532 14044 18596
rect 14108 18532 14109 18596
rect 14043 18531 14109 18532
rect 14046 13837 14106 18531
rect 14043 13836 14109 13837
rect 14043 13772 14044 13836
rect 14108 13772 14109 13836
rect 14043 13771 14109 13772
rect 14230 13701 14290 20843
rect 15518 15197 15578 22611
rect 17723 20772 17789 20773
rect 17723 20708 17724 20772
rect 17788 20708 17789 20772
rect 17723 20707 17789 20708
rect 17355 18052 17421 18053
rect 17355 17988 17356 18052
rect 17420 17988 17421 18052
rect 17355 17987 17421 17988
rect 16251 17508 16317 17509
rect 16251 17444 16252 17508
rect 16316 17444 16317 17508
rect 16251 17443 16317 17444
rect 15515 15196 15581 15197
rect 15515 15132 15516 15196
rect 15580 15132 15581 15196
rect 15515 15131 15581 15132
rect 16254 14653 16314 17443
rect 16251 14652 16317 14653
rect 16251 14588 16252 14652
rect 16316 14588 16317 14652
rect 16251 14587 16317 14588
rect 14227 13700 14293 13701
rect 14227 13636 14228 13700
rect 14292 13636 14293 13700
rect 14227 13635 14293 13636
rect 15147 11252 15213 11253
rect 15147 11188 15148 11252
rect 15212 11188 15213 11252
rect 15147 11187 15213 11188
rect 13675 11116 13741 11117
rect 13675 11052 13676 11116
rect 13740 11052 13741 11116
rect 13675 11051 13741 11052
rect 12939 8396 13005 8397
rect 12939 8332 12940 8396
rect 13004 8332 13005 8396
rect 12939 8331 13005 8332
rect 8339 8260 8405 8261
rect 8339 8196 8340 8260
rect 8404 8196 8405 8260
rect 8339 8195 8405 8196
rect 13491 7172 13557 7173
rect 13491 7108 13492 7172
rect 13556 7108 13557 7172
rect 13491 7107 13557 7108
rect 7235 6492 7301 6493
rect 7235 6428 7236 6492
rect 7300 6428 7301 6492
rect 7235 6427 7301 6428
rect 13494 4861 13554 7107
rect 13678 6221 13738 11051
rect 15150 6493 15210 11187
rect 15331 9484 15397 9485
rect 15331 9420 15332 9484
rect 15396 9420 15397 9484
rect 15331 9419 15397 9420
rect 15147 6492 15213 6493
rect 15147 6428 15148 6492
rect 15212 6428 15213 6492
rect 15147 6427 15213 6428
rect 13675 6220 13741 6221
rect 13675 6156 13676 6220
rect 13740 6156 13741 6220
rect 13675 6155 13741 6156
rect 13491 4860 13557 4861
rect 13491 4796 13492 4860
rect 13556 4796 13557 4860
rect 13491 4795 13557 4796
rect 6683 3636 6749 3637
rect 6683 3572 6684 3636
rect 6748 3572 6749 3636
rect 6683 3571 6749 3572
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 3187 2684 3253 2685
rect 3187 2620 3188 2684
rect 3252 2620 3253 2684
rect 3187 2619 3253 2620
rect 4208 2128 4528 2688
rect 15334 2685 15394 9419
rect 17358 7037 17418 17987
rect 17726 10301 17786 20707
rect 18094 13565 18154 30227
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 20115 17236 20181 17237
rect 20115 17172 20116 17236
rect 20180 17172 20181 17236
rect 20115 17171 20181 17172
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 18091 13564 18157 13565
rect 18091 13500 18092 13564
rect 18156 13500 18157 13564
rect 18091 13499 18157 13500
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 20118 12749 20178 17171
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 20115 12748 20181 12749
rect 20115 12684 20116 12748
rect 20180 12684 20181 12748
rect 20115 12683 20181 12684
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 17723 10300 17789 10301
rect 17723 10236 17724 10300
rect 17788 10236 17789 10300
rect 17723 10235 17789 10236
rect 17726 7581 17786 10235
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19379 9484 19445 9485
rect 19379 9420 19380 9484
rect 19444 9420 19445 9484
rect 19379 9419 19445 9420
rect 19382 8805 19442 9419
rect 19379 8804 19445 8805
rect 19379 8740 19380 8804
rect 19444 8740 19445 8804
rect 19379 8739 19445 8740
rect 19568 8736 19888 9760
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 20299 8940 20365 8941
rect 20299 8876 20300 8940
rect 20364 8876 20365 8940
rect 20299 8875 20365 8876
rect 20115 8804 20181 8805
rect 20115 8740 20116 8804
rect 20180 8740 20181 8804
rect 20115 8739 20181 8740
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19379 8396 19445 8397
rect 19379 8332 19380 8396
rect 19444 8332 19445 8396
rect 19379 8331 19445 8332
rect 17723 7580 17789 7581
rect 17723 7516 17724 7580
rect 17788 7516 17789 7580
rect 17723 7515 17789 7516
rect 17355 7036 17421 7037
rect 17355 6972 17356 7036
rect 17420 6972 17421 7036
rect 17355 6971 17421 6972
rect 19382 6493 19442 8331
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19379 6492 19445 6493
rect 19379 6428 19380 6492
rect 19444 6428 19445 6492
rect 19379 6427 19445 6428
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 20118 4317 20178 8739
rect 20115 4316 20181 4317
rect 20115 4252 20116 4316
rect 20180 4252 20181 4316
rect 20115 4251 20181 4252
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 15331 2684 15397 2685
rect 15331 2620 15332 2684
rect 15396 2620 15397 2684
rect 15331 2619 15397 2620
rect 19568 2208 19888 3232
rect 20302 2957 20362 8875
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 20299 2956 20365 2957
rect 20299 2892 20300 2956
rect 20364 2892 20365 2956
rect 20299 2891 20365 2892
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 24840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 2760 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 26312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1667941163
transform 1 0 8740 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1667941163
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1667941163
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1667941163
transform 1 0 24656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1667941163
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71
timestamp 1667941163
transform 1 0 7636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_147
timestamp 1667941163
transform 1 0 14628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1667941163
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_158
timestamp 1667941163
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1667941163
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1667941163
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1667941163
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1667941163
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_322 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1667941163
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_350
timestamp 1667941163
transform 1 0 33304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1667941163
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_17
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1667941163
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1667941163
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1667941163
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_64
timestamp 1667941163
transform 1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1667941163
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1667941163
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1667941163
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_92
timestamp 1667941163
transform 1 0 9568 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1667941163
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1667941163
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1667941163
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1667941163
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1667941163
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1667941163
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_183
timestamp 1667941163
transform 1 0 17940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_190
timestamp 1667941163
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1667941163
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1667941163
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_211
timestamp 1667941163
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1667941163
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1667941163
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1667941163
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_251
timestamp 1667941163
transform 1 0 24196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_260
timestamp 1667941163
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_267
timestamp 1667941163
transform 1 0 25668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1667941163
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1667941163
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_13
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1667941163
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1667941163
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1667941163
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1667941163
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1667941163
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1667941163
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1667941163
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_127
timestamp 1667941163
transform 1 0 12788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1667941163
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1667941163
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_173
timestamp 1667941163
transform 1 0 17020 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_179
timestamp 1667941163
transform 1 0 17572 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_216
timestamp 1667941163
transform 1 0 20976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_223
timestamp 1667941163
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_237
timestamp 1667941163
transform 1 0 22908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1667941163
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1667941163
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_272
timestamp 1667941163
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_279
timestamp 1667941163
transform 1 0 26772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1667941163
transform 1 0 27416 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_293
timestamp 1667941163
transform 1 0 28060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1667941163
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_9
timestamp 1667941163
transform 1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_18
timestamp 1667941163
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_42
timestamp 1667941163
transform 1 0 4968 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_50
timestamp 1667941163
transform 1 0 5704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_80
timestamp 1667941163
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_88
timestamp 1667941163
transform 1 0 9200 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1667941163
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1667941163
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1667941163
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_187
timestamp 1667941163
transform 1 0 18308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1667941163
transform 1 0 19044 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1667941163
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1667941163
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1667941163
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1667941163
transform 1 0 24840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1667941163
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1667941163
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_298
timestamp 1667941163
transform 1 0 28520 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_310
timestamp 1667941163
transform 1 0 29624 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_322
timestamp 1667941163
transform 1 0 30728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1667941163
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1667941163
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1667941163
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1667941163
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_62
timestamp 1667941163
transform 1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1667941163
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1667941163
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1667941163
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_129
timestamp 1667941163
transform 1 0 12972 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1667941163
transform 1 0 16100 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_184
timestamp 1667941163
transform 1 0 18032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1667941163
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1667941163
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1667941163
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1667941163
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1667941163
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_242
timestamp 1667941163
transform 1 0 23368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1667941163
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_258
timestamp 1667941163
transform 1 0 24840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_266
timestamp 1667941163
transform 1 0 25576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_272
timestamp 1667941163
transform 1 0 26128 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_276
timestamp 1667941163
transform 1 0 26496 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1667941163
transform 1 0 27600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_292
timestamp 1667941163
transform 1 0 27968 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_296
timestamp 1667941163
transform 1 0 28336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_325
timestamp 1667941163
transform 1 0 31004 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_332
timestamp 1667941163
transform 1 0 31648 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_344
timestamp 1667941163
transform 1 0 32752 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1667941163
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1667941163
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1667941163
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1667941163
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1667941163
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1667941163
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_150
timestamp 1667941163
transform 1 0 14904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_156
timestamp 1667941163
transform 1 0 15456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1667941163
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_183
timestamp 1667941163
transform 1 0 17940 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_196
timestamp 1667941163
transform 1 0 19136 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_200
timestamp 1667941163
transform 1 0 19504 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_210
timestamp 1667941163
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_216
timestamp 1667941163
transform 1 0 20976 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1667941163
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_230
timestamp 1667941163
transform 1 0 22264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1667941163
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1667941163
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_258
timestamp 1667941163
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_265
timestamp 1667941163
transform 1 0 25484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1667941163
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_61
timestamp 1667941163
transform 1 0 6716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_98
timestamp 1667941163
transform 1 0 10120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp 1667941163
transform 1 0 10764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1667941163
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp 1667941163
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_171
timestamp 1667941163
transform 1 0 16836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_175
timestamp 1667941163
transform 1 0 17204 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1667941163
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_214
timestamp 1667941163
transform 1 0 20792 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_228
timestamp 1667941163
transform 1 0 22080 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1667941163
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_242
timestamp 1667941163
transform 1 0 23368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1667941163
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_256
timestamp 1667941163
transform 1 0 24656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_260
timestamp 1667941163
transform 1 0 25024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1667941163
transform 1 0 26220 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_278
timestamp 1667941163
transform 1 0 26680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_290
timestamp 1667941163
transform 1 0 27784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1667941163
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_10
timestamp 1667941163
transform 1 0 2024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1667941163
transform 1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1667941163
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1667941163
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1667941163
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1667941163
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_135
timestamp 1667941163
transform 1 0 13524 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_139
timestamp 1667941163
transform 1 0 13892 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1667941163
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1667941163
transform 1 0 18308 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_194
timestamp 1667941163
transform 1 0 18952 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1667941163
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1667941163
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_230
timestamp 1667941163
transform 1 0 22264 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1667941163
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_251
timestamp 1667941163
transform 1 0 24196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_258
timestamp 1667941163
transform 1 0 24840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_262
timestamp 1667941163
transform 1 0 25208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_266
timestamp 1667941163
transform 1 0 25576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_286
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_298
timestamp 1667941163
transform 1 0 28520 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_310
timestamp 1667941163
transform 1 0 29624 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_322
timestamp 1667941163
transform 1 0 30728 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1667941163
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_342
timestamp 1667941163
transform 1 0 32568 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_354
timestamp 1667941163
transform 1 0 33672 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_366
timestamp 1667941163
transform 1 0 34776 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_378
timestamp 1667941163
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1667941163
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_401
timestamp 1667941163
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1667941163
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_33
timestamp 1667941163
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_45
timestamp 1667941163
transform 1 0 5244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_51
timestamp 1667941163
transform 1 0 5796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_72
timestamp 1667941163
transform 1 0 7728 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_78
timestamp 1667941163
transform 1 0 8280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_89
timestamp 1667941163
transform 1 0 9292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1667941163
transform 1 0 9660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1667941163
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1667941163
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1667941163
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_159
timestamp 1667941163
transform 1 0 15732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1667941163
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_183
timestamp 1667941163
transform 1 0 17940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1667941163
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_208
timestamp 1667941163
transform 1 0 20240 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_216
timestamp 1667941163
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_226
timestamp 1667941163
transform 1 0 21896 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_241
timestamp 1667941163
transform 1 0 23276 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_258
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_270
timestamp 1667941163
transform 1 0 25944 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_282
timestamp 1667941163
transform 1 0 27048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_294
timestamp 1667941163
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1667941163
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1667941163
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1667941163
transform 1 0 4048 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_36
timestamp 1667941163
transform 1 0 4416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1667941163
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_47
timestamp 1667941163
transform 1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_70
timestamp 1667941163
transform 1 0 7544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1667941163
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1667941163
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1667941163
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_148
timestamp 1667941163
transform 1 0 14720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_188
timestamp 1667941163
transform 1 0 18400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_196
timestamp 1667941163
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1667941163
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_210
timestamp 1667941163
transform 1 0 20424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1667941163
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1667941163
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1667941163
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_251
timestamp 1667941163
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_256
timestamp 1667941163
transform 1 0 24656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_260
timestamp 1667941163
transform 1 0 25024 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1667941163
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp 1667941163
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_46
timestamp 1667941163
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1667941163
transform 1 0 5704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_72
timestamp 1667941163
transform 1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_78
timestamp 1667941163
transform 1 0 8280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1667941163
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1667941163
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_156
timestamp 1667941163
transform 1 0 15456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1667941163
transform 1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1667941163
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1667941163
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_203
timestamp 1667941163
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_207
timestamp 1667941163
transform 1 0 20148 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_217
timestamp 1667941163
transform 1 0 21068 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1667941163
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_237
timestamp 1667941163
transform 1 0 22908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1667941163
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_270
timestamp 1667941163
transform 1 0 25944 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_282
timestamp 1667941163
transform 1 0 27048 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_294
timestamp 1667941163
transform 1 0 28152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_327
timestamp 1667941163
transform 1 0 31188 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_331
timestamp 1667941163
transform 1 0 31556 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_343
timestamp 1667941163
transform 1 0 32660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1667941163
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_373
timestamp 1667941163
transform 1 0 35420 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1667941163
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_34
timestamp 1667941163
transform 1 0 4232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 1667941163
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_47
timestamp 1667941163
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_62
timestamp 1667941163
transform 1 0 6808 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_68
timestamp 1667941163
transform 1 0 7360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1667941163
transform 1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_96
timestamp 1667941163
transform 1 0 9936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1667941163
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1667941163
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1667941163
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 1667941163
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1667941163
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1667941163
transform 1 0 17572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_196
timestamp 1667941163
transform 1 0 19136 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1667941163
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1667941163
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_230
timestamp 1667941163
transform 1 0 22264 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_246
timestamp 1667941163
transform 1 0 23736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_253
timestamp 1667941163
transform 1 0 24380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_259
timestamp 1667941163
transform 1 0 24932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_263
timestamp 1667941163
transform 1 0 25300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp 1667941163
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1667941163
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_345
timestamp 1667941163
transform 1 0 32844 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_401
timestamp 1667941163
transform 1 0 37996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1667941163
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_42
timestamp 1667941163
transform 1 0 4968 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_51
timestamp 1667941163
transform 1 0 5796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1667941163
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1667941163
transform 1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1667941163
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_123
timestamp 1667941163
transform 1 0 12420 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_131
timestamp 1667941163
transform 1 0 13156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_163
timestamp 1667941163
transform 1 0 16100 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_179
timestamp 1667941163
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1667941163
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_208
timestamp 1667941163
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1667941163
transform 1 0 20884 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1667941163
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_235
timestamp 1667941163
transform 1 0 22724 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_242
timestamp 1667941163
transform 1 0 23368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1667941163
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_314
timestamp 1667941163
transform 1 0 29992 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_326
timestamp 1667941163
transform 1 0 31096 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_338
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_350
timestamp 1667941163
transform 1 0 33304 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1667941163
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_25
timestamp 1667941163
transform 1 0 3404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_33
timestamp 1667941163
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_62
timestamp 1667941163
transform 1 0 6808 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_68
timestamp 1667941163
transform 1 0 7360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_92
timestamp 1667941163
transform 1 0 9568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1667941163
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1667941163
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1667941163
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_159
timestamp 1667941163
transform 1 0 15732 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_180
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_197
timestamp 1667941163
transform 1 0 19228 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_207
timestamp 1667941163
transform 1 0 20148 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_213
timestamp 1667941163
transform 1 0 20700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1667941163
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_244
timestamp 1667941163
transform 1 0 23552 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_252
timestamp 1667941163
transform 1 0 24288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_262
timestamp 1667941163
transform 1 0 25208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1667941163
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1667941163
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_54
timestamp 1667941163
transform 1 0 6072 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_107
timestamp 1667941163
transform 1 0 10948 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_115
timestamp 1667941163
transform 1 0 11684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1667941163
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1667941163
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_171
timestamp 1667941163
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_184
timestamp 1667941163
transform 1 0 18032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_208
timestamp 1667941163
transform 1 0 20240 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_216
timestamp 1667941163
transform 1 0 20976 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_226
timestamp 1667941163
transform 1 0 21896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1667941163
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_238
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1667941163
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_272
timestamp 1667941163
transform 1 0 26128 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_284
timestamp 1667941163
transform 1 0 27232 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_296
timestamp 1667941163
transform 1 0 28336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_16
timestamp 1667941163
transform 1 0 2576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1667941163
transform 1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1667941163
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1667941163
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_94
timestamp 1667941163
transform 1 0 9752 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1667941163
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_136
timestamp 1667941163
transform 1 0 13616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1667941163
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_179
timestamp 1667941163
transform 1 0 17572 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_200
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1667941163
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_239
timestamp 1667941163
transform 1 0 23092 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_246
timestamp 1667941163
transform 1 0 23736 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_253
timestamp 1667941163
transform 1 0 24380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_260
timestamp 1667941163
transform 1 0 25024 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1667941163
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_309
timestamp 1667941163
transform 1 0 29532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_321
timestamp 1667941163
transform 1 0 30636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1667941163
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1667941163
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1667941163
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1667941163
transform 1 0 6256 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1667941163
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_91
timestamp 1667941163
transform 1 0 9476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_98
timestamp 1667941163
transform 1 0 10120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_105
timestamp 1667941163
transform 1 0 10764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_129
timestamp 1667941163
transform 1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1667941163
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1667941163
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1667941163
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1667941163
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_223
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1667941163
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1667941163
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_258
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_273
timestamp 1667941163
transform 1 0 26220 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_280
timestamp 1667941163
transform 1 0 26864 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_292
timestamp 1667941163
transform 1 0 27968 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1667941163
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_28
timestamp 1667941163
transform 1 0 3680 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_63
timestamp 1667941163
transform 1 0 6900 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_70
timestamp 1667941163
transform 1 0 7544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_95
timestamp 1667941163
transform 1 0 9844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1667941163
transform 1 0 10212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1667941163
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1667941163
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1667941163
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_180
timestamp 1667941163
transform 1 0 17664 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1667941163
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_202
timestamp 1667941163
transform 1 0 19688 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_208
timestamp 1667941163
transform 1 0 20240 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_240
timestamp 1667941163
transform 1 0 23184 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_248
timestamp 1667941163
transform 1 0 23920 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_253
timestamp 1667941163
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1667941163
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_264
timestamp 1667941163
transform 1 0 25392 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_268
timestamp 1667941163
transform 1 0 25760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_309
timestamp 1667941163
transform 1 0 29532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_313
timestamp 1667941163
transform 1 0 29900 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1667941163
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1667941163
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1667941163
transform 1 0 5796 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1667941163
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1667941163
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1667941163
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_106
timestamp 1667941163
transform 1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_131
timestamp 1667941163
transform 1 0 13156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1667941163
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1667941163
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_205
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_222
timestamp 1667941163
transform 1 0 21528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_236
timestamp 1667941163
transform 1 0 22816 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_243
timestamp 1667941163
transform 1 0 23460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1667941163
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_314
timestamp 1667941163
transform 1 0 29992 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_326
timestamp 1667941163
transform 1 0 31096 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_338
timestamp 1667941163
transform 1 0 32200 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_350
timestamp 1667941163
transform 1 0 33304 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1667941163
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_26
timestamp 1667941163
transform 1 0 3496 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1667941163
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1667941163
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1667941163
transform 1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1667941163
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1667941163
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1667941163
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1667941163
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1667941163
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_244
timestamp 1667941163
transform 1 0 23552 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_256
timestamp 1667941163
transform 1 0 24656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_268
timestamp 1667941163
transform 1 0 25760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1667941163
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_42
timestamp 1667941163
transform 1 0 4968 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_50
timestamp 1667941163
transform 1 0 5704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_71
timestamp 1667941163
transform 1 0 7636 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1667941163
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1667941163
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1667941163
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1667941163
transform 1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_180
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1667941163
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1667941163
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1667941163
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1667941163
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_225
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_231
timestamp 1667941163
transform 1 0 22356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_235
timestamp 1667941163
transform 1 0 22724 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_243
timestamp 1667941163
transform 1 0 23460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_271
timestamp 1667941163
transform 1 0 26036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_280
timestamp 1667941163
transform 1 0 26864 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_287
timestamp 1667941163
transform 1 0 27508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_299
timestamp 1667941163
transform 1 0 28612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_25
timestamp 1667941163
transform 1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1667941163
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1667941163
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1667941163
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1667941163
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_152
timestamp 1667941163
transform 1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_156
timestamp 1667941163
transform 1 0 15456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1667941163
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1667941163
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_229
timestamp 1667941163
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1667941163
transform 1 0 23000 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_245
timestamp 1667941163
transform 1 0 23644 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_257
timestamp 1667941163
transform 1 0 24748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_269
timestamp 1667941163
transform 1 0 25852 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1667941163
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_353
timestamp 1667941163
transform 1 0 33580 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_357
timestamp 1667941163
transform 1 0 33948 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_369
timestamp 1667941163
transform 1 0 35052 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_381
timestamp 1667941163
transform 1 0 36156 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_389
timestamp 1667941163
transform 1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1667941163
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_36
timestamp 1667941163
transform 1 0 4416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1667941163
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1667941163
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_75
timestamp 1667941163
transform 1 0 8004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1667941163
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1667941163
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1667941163
transform 1 0 14812 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_168
timestamp 1667941163
transform 1 0 16560 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_185
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_207
timestamp 1667941163
transform 1 0 20148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_214
timestamp 1667941163
transform 1 0 20792 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_222
timestamp 1667941163
transform 1 0 21528 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_227
timestamp 1667941163
transform 1 0 21988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1667941163
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_263
timestamp 1667941163
transform 1 0 25300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_275
timestamp 1667941163
transform 1 0 26404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1667941163
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_295
timestamp 1667941163
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_371
timestamp 1667941163
transform 1 0 35236 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_375
timestamp 1667941163
transform 1 0 35604 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_387
timestamp 1667941163
transform 1 0 36708 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_399
timestamp 1667941163
transform 1 0 37812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_25
timestamp 1667941163
transform 1 0 3404 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_64
timestamp 1667941163
transform 1 0 6992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1667941163
transform 1 0 7636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_98
timestamp 1667941163
transform 1 0 10120 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_106
timestamp 1667941163
transform 1 0 10856 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1667941163
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_153
timestamp 1667941163
transform 1 0 15180 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_191
timestamp 1667941163
transform 1 0 18676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_242
timestamp 1667941163
transform 1 0 23368 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_248
timestamp 1667941163
transform 1 0 23920 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_252
timestamp 1667941163
transform 1 0 24288 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_264
timestamp 1667941163
transform 1 0 25392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1667941163
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_291
timestamp 1667941163
transform 1 0 27876 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_302
timestamp 1667941163
transform 1 0 28888 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_314
timestamp 1667941163
transform 1 0 29992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1667941163
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1667941163
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_402
timestamp 1667941163
transform 1 0 38088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1667941163
transform 1 0 38456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1667941163
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1667941163
transform 1 0 5796 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1667941163
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_89
timestamp 1667941163
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1667941163
transform 1 0 9660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_117
timestamp 1667941163
transform 1 0 11868 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1667941163
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_166
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_174
timestamp 1667941163
transform 1 0 17112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1667941163
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1667941163
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_208
timestamp 1667941163
transform 1 0 20240 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_216
timestamp 1667941163
transform 1 0 20976 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1667941163
transform 1 0 23184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_263
timestamp 1667941163
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_275
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_287
timestamp 1667941163
transform 1 0 27508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_295
timestamp 1667941163
transform 1 0 28244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_88
timestamp 1667941163
transform 1 0 9200 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_94
timestamp 1667941163
transform 1 0 9752 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1667941163
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1667941163
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1667941163
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_157
timestamp 1667941163
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_180
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1667941163
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_210
timestamp 1667941163
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1667941163
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_240
timestamp 1667941163
transform 1 0 23184 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_248
timestamp 1667941163
transform 1 0 23920 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_254
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_266
timestamp 1667941163
transform 1 0 25576 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_272
timestamp 1667941163
transform 1 0 26128 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1667941163
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_291
timestamp 1667941163
transform 1 0 27876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1667941163
transform 1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_42
timestamp 1667941163
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_46
timestamp 1667941163
transform 1 0 5336 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1667941163
transform 1 0 7268 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_91
timestamp 1667941163
transform 1 0 9476 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_98
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_105
timestamp 1667941163
transform 1 0 10764 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_129
timestamp 1667941163
transform 1 0 12972 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_147
timestamp 1667941163
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_154
timestamp 1667941163
transform 1 0 15272 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_160
timestamp 1667941163
transform 1 0 15824 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1667941163
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1667941163
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1667941163
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1667941163
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1667941163
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_211
timestamp 1667941163
transform 1 0 20516 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_215
timestamp 1667941163
transform 1 0 20884 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_227
timestamp 1667941163
transform 1 0 21988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_242
timestamp 1667941163
transform 1 0 23368 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_246
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1667941163
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_268
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_280
timestamp 1667941163
transform 1 0 26864 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_288
timestamp 1667941163
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_293
timestamp 1667941163
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1667941163
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_28
timestamp 1667941163
transform 1 0 3680 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_63
timestamp 1667941163
transform 1 0 6900 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_71
timestamp 1667941163
transform 1 0 7636 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1667941163
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_138
timestamp 1667941163
transform 1 0 13800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1667941163
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_185
timestamp 1667941163
transform 1 0 18124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_197
timestamp 1667941163
transform 1 0 19228 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_205
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_209
timestamp 1667941163
transform 1 0 20332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1667941163
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_246
timestamp 1667941163
transform 1 0 23736 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_265
timestamp 1667941163
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1667941163
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_357
timestamp 1667941163
transform 1 0 33948 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_363
timestamp 1667941163
transform 1 0 34500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_375
timestamp 1667941163
transform 1 0 35604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_387
timestamp 1667941163
transform 1 0 36708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_61
timestamp 1667941163
transform 1 0 6716 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1667941163
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 1667941163
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1667941163
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1667941163
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1667941163
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1667941163
transform 1 0 20424 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_222
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_25
timestamp 1667941163
transform 1 0 3404 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1667941163
transform 1 0 3956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1667941163
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1667941163
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1667941163
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_136
timestamp 1667941163
transform 1 0 13616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_153
timestamp 1667941163
transform 1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1667941163
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_187
timestamp 1667941163
transform 1 0 18308 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_207
timestamp 1667941163
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_243
timestamp 1667941163
transform 1 0 23460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_250
timestamp 1667941163
transform 1 0 24104 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1667941163
transform 1 0 24840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1667941163
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1667941163
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_369
timestamp 1667941163
transform 1 0 35052 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_92
timestamp 1667941163
transform 1 0 9568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1667941163
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_116
timestamp 1667941163
transform 1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_123
timestamp 1667941163
transform 1 0 12420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_131
timestamp 1667941163
transform 1 0 13156 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1667941163
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_159
timestamp 1667941163
transform 1 0 15732 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1667941163
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1667941163
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_211
timestamp 1667941163
transform 1 0 20516 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_223
timestamp 1667941163
transform 1 0 21620 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_235
timestamp 1667941163
transform 1 0 22724 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_267
timestamp 1667941163
transform 1 0 25668 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_274
timestamp 1667941163
transform 1 0 26312 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_286
timestamp 1667941163
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1667941163
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1667941163
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1667941163
transform 1 0 2760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_26
timestamp 1667941163
transform 1 0 3496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_30
timestamp 1667941163
transform 1 0 3864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_64
timestamp 1667941163
transform 1 0 6992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_88
timestamp 1667941163
transform 1 0 9200 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1667941163
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_135
timestamp 1667941163
transform 1 0 13524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1667941163
transform 1 0 15272 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_174
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_180
timestamp 1667941163
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_194
timestamp 1667941163
transform 1 0 18952 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_202
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_209
timestamp 1667941163
transform 1 0 20332 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_238
timestamp 1667941163
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_243
timestamp 1667941163
transform 1 0 23460 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_250
timestamp 1667941163
transform 1 0 24104 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_256
timestamp 1667941163
transform 1 0 24656 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 1667941163
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1667941163
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_316
timestamp 1667941163
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1667941163
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_401
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1667941163
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_38
timestamp 1667941163
transform 1 0 4600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_55
timestamp 1667941163
transform 1 0 6164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1667941163
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_131
timestamp 1667941163
transform 1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_156
timestamp 1667941163
transform 1 0 15456 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_164
timestamp 1667941163
transform 1 0 16192 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1667941163
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 1667941163
transform 1 0 16928 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_176
timestamp 1667941163
transform 1 0 17296 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1667941163
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_217
timestamp 1667941163
transform 1 0 21068 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_229
timestamp 1667941163
transform 1 0 22172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1667941163
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_240
timestamp 1667941163
transform 1 0 23184 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_258
timestamp 1667941163
transform 1 0 24840 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_266
timestamp 1667941163
transform 1 0 25576 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_271
timestamp 1667941163
transform 1 0 26036 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_283
timestamp 1667941163
transform 1 0 27140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_295
timestamp 1667941163
transform 1 0 28244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_339
timestamp 1667941163
transform 1 0 32292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_351
timestamp 1667941163
transform 1 0 33396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_18
timestamp 1667941163
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_31
timestamp 1667941163
transform 1 0 3956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_44
timestamp 1667941163
transform 1 0 5152 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_50
timestamp 1667941163
transform 1 0 5704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_68
timestamp 1667941163
transform 1 0 7360 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_74
timestamp 1667941163
transform 1 0 7912 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_88
timestamp 1667941163
transform 1 0 9200 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_97
timestamp 1667941163
transform 1 0 10028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_128
timestamp 1667941163
transform 1 0 12880 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_136
timestamp 1667941163
transform 1 0 13616 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_150
timestamp 1667941163
transform 1 0 14904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1667941163
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1667941163
transform 1 0 17664 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_186
timestamp 1667941163
transform 1 0 18216 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_200
timestamp 1667941163
transform 1 0 19504 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_212
timestamp 1667941163
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1667941163
transform 1 0 23460 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_247
timestamp 1667941163
transform 1 0 23828 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_254
timestamp 1667941163
transform 1 0 24472 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1667941163
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_34
timestamp 1667941163
transform 1 0 4232 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1667941163
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_60
timestamp 1667941163
transform 1 0 6624 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1667941163
transform 1 0 9568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_115
timestamp 1667941163
transform 1 0 11684 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_119
timestamp 1667941163
transform 1 0 12052 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1667941163
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1667941163
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_159
timestamp 1667941163
transform 1 0 15732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_166
timestamp 1667941163
transform 1 0 16376 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_183
timestamp 1667941163
transform 1 0 17940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_213
timestamp 1667941163
transform 1 0 20700 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_225
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_237
timestamp 1667941163
transform 1 0 22908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_257
timestamp 1667941163
transform 1 0 24748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_261
timestamp 1667941163
transform 1 0 25116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_268
timestamp 1667941163
transform 1 0 25760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_275
timestamp 1667941163
transform 1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_282
timestamp 1667941163
transform 1 0 27048 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_294
timestamp 1667941163
transform 1 0 28152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_326
timestamp 1667941163
transform 1 0 31096 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_338
timestamp 1667941163
transform 1 0 32200 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_19
timestamp 1667941163
transform 1 0 2852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_32
timestamp 1667941163
transform 1 0 4048 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_78
timestamp 1667941163
transform 1 0 8280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_91
timestamp 1667941163
transform 1 0 9476 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_99
timestamp 1667941163
transform 1 0 10212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1667941163
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1667941163
transform 1 0 12788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_140
timestamp 1667941163
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_152
timestamp 1667941163
transform 1 0 15088 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_160
timestamp 1667941163
transform 1 0 15824 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1667941163
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_187
timestamp 1667941163
transform 1 0 18308 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1667941163
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_198
timestamp 1667941163
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_211
timestamp 1667941163
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_235
timestamp 1667941163
transform 1 0 22724 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_247
timestamp 1667941163
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_259
timestamp 1667941163
transform 1 0 24932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_264
timestamp 1667941163
transform 1 0 25392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_268
timestamp 1667941163
transform 1 0 25760 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_342
timestamp 1667941163
transform 1 0 32568 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_354
timestamp 1667941163
transform 1 0 33672 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_366
timestamp 1667941163
transform 1 0 34776 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_378
timestamp 1667941163
transform 1 0 35880 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1667941163
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1667941163
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 1667941163
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_37
timestamp 1667941163
transform 1 0 4508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_44
timestamp 1667941163
transform 1 0 5152 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp 1667941163
transform 1 0 5796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_58
timestamp 1667941163
transform 1 0 6440 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_64
timestamp 1667941163
transform 1 0 6992 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_68
timestamp 1667941163
transform 1 0 7360 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1667941163
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1667941163
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_113
timestamp 1667941163
transform 1 0 11500 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1667941163
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_131
timestamp 1667941163
transform 1 0 13156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_147
timestamp 1667941163
transform 1 0 14628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_164
timestamp 1667941163
transform 1 0 16192 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_181
timestamp 1667941163
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_214
timestamp 1667941163
transform 1 0 20792 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_222
timestamp 1667941163
transform 1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_227
timestamp 1667941163
transform 1 0 21988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_239
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_261
timestamp 1667941163
transform 1 0 25116 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_275
timestamp 1667941163
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1667941163
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1667941163
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_402
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1667941163
transform 1 0 38456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1667941163
transform 1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_29
timestamp 1667941163
transform 1 0 3772 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_36
timestamp 1667941163
transform 1 0 4416 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_42
timestamp 1667941163
transform 1 0 4968 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_46
timestamp 1667941163
transform 1 0 5336 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_50
timestamp 1667941163
transform 1 0 5704 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1667941163
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_65
timestamp 1667941163
transform 1 0 7084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_72
timestamp 1667941163
transform 1 0 7728 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_80
timestamp 1667941163
transform 1 0 8464 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_85
timestamp 1667941163
transform 1 0 8924 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_92
timestamp 1667941163
transform 1 0 9568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1667941163
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_122
timestamp 1667941163
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1667941163
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_153
timestamp 1667941163
transform 1 0 15180 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_158
timestamp 1667941163
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1667941163
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_188
timestamp 1667941163
transform 1 0 18400 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_200
timestamp 1667941163
transform 1 0 19504 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_212
timestamp 1667941163
transform 1 0 20608 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1667941163
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1667941163
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1667941163
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_39
timestamp 1667941163
transform 1 0 4692 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_43
timestamp 1667941163
transform 1 0 5060 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_54
timestamp 1667941163
transform 1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_61
timestamp 1667941163
transform 1 0 6716 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_68
timestamp 1667941163
transform 1 0 7360 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1667941163
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_104
timestamp 1667941163
transform 1 0 10672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_117
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_125
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_146
timestamp 1667941163
transform 1 0 14536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_150
timestamp 1667941163
transform 1 0 14904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_160
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_185
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1667941163
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_208
timestamp 1667941163
transform 1 0 20240 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_220
timestamp 1667941163
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_232
timestamp 1667941163
transform 1 0 22448 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_242
timestamp 1667941163
transform 1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_317
timestamp 1667941163
transform 1 0 30268 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_322
timestamp 1667941163
transform 1 0 30728 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_334
timestamp 1667941163
transform 1 0 31832 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_346
timestamp 1667941163
transform 1 0 32936 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_358
timestamp 1667941163
transform 1 0 34040 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_12
timestamp 1667941163
transform 1 0 2208 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_20
timestamp 1667941163
transform 1 0 2944 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_31
timestamp 1667941163
transform 1 0 3956 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_38
timestamp 1667941163
transform 1 0 4600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_45
timestamp 1667941163
transform 1 0 5244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1667941163
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_76
timestamp 1667941163
transform 1 0 8096 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_89
timestamp 1667941163
transform 1 0 9292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_96
timestamp 1667941163
transform 1 0 9936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_103
timestamp 1667941163
transform 1 0 10580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_119
timestamp 1667941163
transform 1 0 12052 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_132
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1667941163
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_152
timestamp 1667941163
transform 1 0 15088 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_160
timestamp 1667941163
transform 1 0 15824 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1667941163
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_186
timestamp 1667941163
transform 1 0 18216 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_194
timestamp 1667941163
transform 1 0 18952 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_203
timestamp 1667941163
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1667941163
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1667941163
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_240
timestamp 1667941163
transform 1 0 23184 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_244
timestamp 1667941163
transform 1 0 23552 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_256
timestamp 1667941163
transform 1 0 24656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_268
timestamp 1667941163
transform 1 0 25760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_325
timestamp 1667941163
transform 1 0 31004 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1667941163
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1667941163
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1667941163
transform 1 0 2116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_18
timestamp 1667941163
transform 1 0 2760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1667941163
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_36
timestamp 1667941163
transform 1 0 4416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_43
timestamp 1667941163
transform 1 0 5060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_50
timestamp 1667941163
transform 1 0 5704 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_57
timestamp 1667941163
transform 1 0 6348 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_63
timestamp 1667941163
transform 1 0 6900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_67
timestamp 1667941163
transform 1 0 7268 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1667941163
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1667941163
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_105
timestamp 1667941163
transform 1 0 10764 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_112
timestamp 1667941163
transform 1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_120
timestamp 1667941163
transform 1 0 12144 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1667941163
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1667941163
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_174
timestamp 1667941163
transform 1 0 17112 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_182
timestamp 1667941163
transform 1 0 17848 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1667941163
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_202
timestamp 1667941163
transform 1 0 19688 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_217
timestamp 1667941163
transform 1 0 21068 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_229
timestamp 1667941163
transform 1 0 22172 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_235
timestamp 1667941163
transform 1 0 22724 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_239
timestamp 1667941163
transform 1 0 23092 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_243
timestamp 1667941163
transform 1 0 23460 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1667941163
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_13
timestamp 1667941163
transform 1 0 2300 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_28
timestamp 1667941163
transform 1 0 3680 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_32
timestamp 1667941163
transform 1 0 4048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_46
timestamp 1667941163
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_73
timestamp 1667941163
transform 1 0 7820 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_83
timestamp 1667941163
transform 1 0 8740 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_96
timestamp 1667941163
transform 1 0 9936 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1667941163
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_119
timestamp 1667941163
transform 1 0 12052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1667941163
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_148
timestamp 1667941163
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_155
timestamp 1667941163
transform 1 0 15364 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1667941163
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_192
timestamp 1667941163
transform 1 0 18768 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_204
timestamp 1667941163
transform 1 0 19872 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_213
timestamp 1667941163
transform 1 0 20700 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1667941163
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_236
timestamp 1667941163
transform 1 0 22816 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1667941163
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_254
timestamp 1667941163
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_266
timestamp 1667941163
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1667941163
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_301
timestamp 1667941163
transform 1 0 28796 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_306
timestamp 1667941163
transform 1 0 29256 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_318
timestamp 1667941163
transform 1 0 30360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1667941163
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_22
timestamp 1667941163
transform 1 0 3128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_34
timestamp 1667941163
transform 1 0 4232 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_48
timestamp 1667941163
transform 1 0 5520 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 1667941163
transform 1 0 6624 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1667941163
transform 1 0 9476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_95
timestamp 1667941163
transform 1 0 9844 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_104
timestamp 1667941163
transform 1 0 10672 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_119
timestamp 1667941163
transform 1 0 12052 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_131
timestamp 1667941163
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_169
timestamp 1667941163
transform 1 0 16652 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1667941163
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_203
timestamp 1667941163
transform 1 0 19780 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_211
timestamp 1667941163
transform 1 0 20516 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_216
timestamp 1667941163
transform 1 0 20976 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_228
timestamp 1667941163
transform 1 0 22080 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_240
timestamp 1667941163
transform 1 0 23184 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_283
timestamp 1667941163
transform 1 0 27140 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_287
timestamp 1667941163
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1667941163
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_337
timestamp 1667941163
transform 1 0 32108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_341
timestamp 1667941163
transform 1 0 32476 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_353
timestamp 1667941163
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1667941163
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_14
timestamp 1667941163
transform 1 0 2392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_21
timestamp 1667941163
transform 1 0 3036 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_28
timestamp 1667941163
transform 1 0 3680 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_35
timestamp 1667941163
transform 1 0 4324 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_42
timestamp 1667941163
transform 1 0 4968 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1667941163
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_89
timestamp 1667941163
transform 1 0 9292 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1667941163
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_121
timestamp 1667941163
transform 1 0 12236 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_126
timestamp 1667941163
transform 1 0 12696 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_138
timestamp 1667941163
transform 1 0 13800 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_144
timestamp 1667941163
transform 1 0 14352 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_156
timestamp 1667941163
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_174
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_182
timestamp 1667941163
transform 1 0 17848 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_186
timestamp 1667941163
transform 1 0 18216 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_194
timestamp 1667941163
transform 1 0 18952 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_201
timestamp 1667941163
transform 1 0 19596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1667941163
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1667941163
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_13
timestamp 1667941163
transform 1 0 2300 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1667941163
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_34
timestamp 1667941163
transform 1 0 4232 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_46
timestamp 1667941163
transform 1 0 5336 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_54
timestamp 1667941163
transform 1 0 6072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_59
timestamp 1667941163
transform 1 0 6532 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_66
timestamp 1667941163
transform 1 0 7176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_78
timestamp 1667941163
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_93
timestamp 1667941163
transform 1 0 9660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_103
timestamp 1667941163
transform 1 0 10580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_115
timestamp 1667941163
transform 1 0 11684 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_122
timestamp 1667941163
transform 1 0 12328 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1667941163
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_156
timestamp 1667941163
transform 1 0 15456 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_160
timestamp 1667941163
transform 1 0 15824 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_174
timestamp 1667941163
transform 1 0 17112 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_182
timestamp 1667941163
transform 1 0 17848 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1667941163
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_202
timestamp 1667941163
transform 1 0 19688 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_217
timestamp 1667941163
transform 1 0 21068 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_232
timestamp 1667941163
transform 1 0 22448 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_239
timestamp 1667941163
transform 1 0 23092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_7
timestamp 1667941163
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1667941163
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_18
timestamp 1667941163
transform 1 0 2760 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_25
timestamp 1667941163
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_37
timestamp 1667941163
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_49
timestamp 1667941163
transform 1 0 5612 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_64
timestamp 1667941163
transform 1 0 6992 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_72
timestamp 1667941163
transform 1 0 7728 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1667941163
transform 1 0 8188 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_90
timestamp 1667941163
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_102
timestamp 1667941163
transform 1 0 10488 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1667941163
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp 1667941163
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_141
timestamp 1667941163
transform 1 0 14076 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_148
timestamp 1667941163
transform 1 0 14720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1667941163
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_342
timestamp 1667941163
transform 1 0 32568 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_354
timestamp 1667941163
transform 1 0 33672 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_366
timestamp 1667941163
transform 1 0 34776 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_378
timestamp 1667941163
transform 1 0 35880 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1667941163
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_16
timestamp 1667941163
transform 1 0 2576 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_115
timestamp 1667941163
transform 1 0 11684 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1667941163
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_131
timestamp 1667941163
transform 1 0 13156 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_146
timestamp 1667941163
transform 1 0 14536 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_158
timestamp 1667941163
transform 1 0 15640 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_170
timestamp 1667941163
transform 1 0 16744 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_182
timestamp 1667941163
transform 1 0 17848 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_295
timestamp 1667941163
transform 1 0 28244 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1667941163
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1667941163
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1667941163
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1667941163
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_180
timestamp 1667941163
transform 1 0 17664 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_191
timestamp 1667941163
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_203
timestamp 1667941163
transform 1 0 19780 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_215
timestamp 1667941163
transform 1 0 20884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_309
timestamp 1667941163
transform 1 0 29532 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_321
timestamp 1667941163
transform 1 0 30636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_333
timestamp 1667941163
transform 1 0 31740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_342
timestamp 1667941163
transform 1 0 32568 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_354
timestamp 1667941163
transform 1 0 33672 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_366
timestamp 1667941163
transform 1 0 34776 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_378
timestamp 1667941163
transform 1 0 35880 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_390
timestamp 1667941163
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_401
timestamp 1667941163
transform 1 0 37996 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_149
timestamp 1667941163
transform 1 0 14812 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_155
timestamp 1667941163
transform 1 0 15364 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_167
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_179
timestamp 1667941163
transform 1 0 17572 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1667941163
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_276
timestamp 1667941163
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_288
timestamp 1667941163
transform 1 0 27600 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_300
timestamp 1667941163
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_68
timestamp 1667941163
transform 1 0 7360 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_80
timestamp 1667941163
transform 1 0 8464 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_92
timestamp 1667941163
transform 1 0 9568 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1667941163
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_352
timestamp 1667941163
transform 1 0 33488 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_364
timestamp 1667941163
transform 1 0 34592 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_376
timestamp 1667941163
transform 1 0 35696 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1667941163
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_59
timestamp 1667941163
transform 1 0 6532 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_63
timestamp 1667941163
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_75
timestamp 1667941163
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_90
timestamp 1667941163
transform 1 0 9384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_102
timestamp 1667941163
transform 1 0 10488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_114
timestamp 1667941163
transform 1 0 11592 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_126
timestamp 1667941163
transform 1 0 12696 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1667941163
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_9
timestamp 1667941163
transform 1 0 1932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_21
timestamp 1667941163
transform 1 0 3036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_33
timestamp 1667941163
transform 1 0 4140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_45
timestamp 1667941163
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1667941163
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_121
timestamp 1667941163
transform 1 0 12236 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1667941163
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_286
timestamp 1667941163
transform 1 0 27416 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_298
timestamp 1667941163
transform 1 0 28520 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_310
timestamp 1667941163
transform 1 0 29624 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_322
timestamp 1667941163
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1667941163
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_45
timestamp 1667941163
transform 1 0 5244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_57
timestamp 1667941163
transform 1 0 6348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_69
timestamp 1667941163
transform 1 0 7452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1667941163
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_89
timestamp 1667941163
transform 1 0 9292 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_93
timestamp 1667941163
transform 1 0 9660 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_105
timestamp 1667941163
transform 1 0 10764 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_117
timestamp 1667941163
transform 1 0 11868 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_129
timestamp 1667941163
transform 1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 1667941163
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_227
timestamp 1667941163
transform 1 0 21988 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_231
timestamp 1667941163
transform 1 0 22356 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1667941163
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_65
timestamp 1667941163
transform 1 0 7084 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_71
timestamp 1667941163
transform 1 0 7636 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_83
timestamp 1667941163
transform 1 0 8740 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_95
timestamp 1667941163
transform 1 0 9844 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1667941163
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_245
timestamp 1667941163
transform 1 0 23644 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_251
timestamp 1667941163
transform 1 0 24196 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_263
timestamp 1667941163
transform 1 0 25300 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_275
timestamp 1667941163
transform 1 0 26404 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_302
timestamp 1667941163
transform 1 0 28888 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_314
timestamp 1667941163
transform 1 0 29992 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_326
timestamp 1667941163
transform 1 0 31096 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1667941163
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1667941163
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_40
timestamp 1667941163
transform 1 0 4784 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_52
timestamp 1667941163
transform 1 0 5888 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_64
timestamp 1667941163
transform 1 0 6992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_68
timestamp 1667941163
transform 1 0 7360 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_72
timestamp 1667941163
transform 1 0 7728 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_90
timestamp 1667941163
transform 1 0 9384 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_102
timestamp 1667941163
transform 1 0 10488 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_114
timestamp 1667941163
transform 1 0 11592 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_126
timestamp 1667941163
transform 1 0 12696 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_159
timestamp 1667941163
transform 1 0 15732 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_163
timestamp 1667941163
transform 1 0 16100 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_175
timestamp 1667941163
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_187
timestamp 1667941163
transform 1 0 18308 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_227
timestamp 1667941163
transform 1 0 21988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_239
timestamp 1667941163
transform 1 0 23092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_258
timestamp 1667941163
transform 1 0 24840 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_270
timestamp 1667941163
transform 1 0 25944 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_282
timestamp 1667941163
transform 1 0 27048 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_294
timestamp 1667941163
transform 1 0 28152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1667941163
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_85
timestamp 1667941163
transform 1 0 8924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_89
timestamp 1667941163
transform 1 0 9292 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_101
timestamp 1667941163
transform 1 0 10396 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_109
timestamp 1667941163
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_49
timestamp 1667941163
transform 1 0 5612 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1667941163
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1667941163
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1667941163
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1667941163
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1667941163
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_197
timestamp 1667941163
transform 1 0 19228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_209
timestamp 1667941163
transform 1 0 20332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1667941163
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_141
timestamp 1667941163
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_145
timestamp 1667941163
transform 1 0 14444 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_157
timestamp 1667941163
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1667941163
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_369
timestamp 1667941163
transform 1 0 35052 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_374
timestamp 1667941163
transform 1 0 35512 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_381
timestamp 1667941163
transform 1 0 36156 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1667941163
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_8
timestamp 1667941163
transform 1 0 1840 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_20
timestamp 1667941163
transform 1 0 2944 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1667941163
transform 1 0 37720 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1667941163
transform 1 0 38456 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_21
timestamp 1667941163
transform 1 0 3036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_33
timestamp 1667941163
transform 1 0 4140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_45
timestamp 1667941163
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1667941163
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_16
timestamp 1667941163
transform 1 0 2576 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_373
timestamp 1667941163
transform 1 0 35420 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_385
timestamp 1667941163
transform 1 0 36524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_22
timestamp 1667941163
transform 1 0 3128 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_34
timestamp 1667941163
transform 1 0 4232 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_46
timestamp 1667941163
transform 1 0 5336 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_85
timestamp 1667941163
transform 1 0 8924 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_91
timestamp 1667941163
transform 1 0 9476 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_103
timestamp 1667941163
transform 1 0 10580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_134
timestamp 1667941163
transform 1 0 13432 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_142
timestamp 1667941163
transform 1 0 14168 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_146
timestamp 1667941163
transform 1 0 14536 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_158
timestamp 1667941163
transform 1 0 15640 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_175
timestamp 1667941163
transform 1 0 17204 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_187
timestamp 1667941163
transform 1 0 18308 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_199
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_211
timestamp 1667941163
transform 1 0 20516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_231
timestamp 1667941163
transform 1 0 22356 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_239
timestamp 1667941163
transform 1 0 23092 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_251
timestamp 1667941163
transform 1 0 24196 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_263
timestamp 1667941163
transform 1 0 25300 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1667941163
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_369
timestamp 1667941163
transform 1 0 35052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_375
timestamp 1667941163
transform 1 0 35604 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_382
timestamp 1667941163
transform 1 0 36248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_70
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_89
timestamp 1667941163
transform 1 0 9292 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_92
timestamp 1667941163
transform 1 0 9568 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1667941163
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_155
timestamp 1667941163
transform 1 0 15364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_160
timestamp 1667941163
transform 1 0 15824 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_177
timestamp 1667941163
transform 1 0 17388 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_182
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1667941163
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1667941163
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0390_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26128 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0392_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0393_
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0394_
timestamp 1667941163
transform 1 0 26772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0395_
timestamp 1667941163
transform 1 0 25760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0397_
timestamp 1667941163
transform 1 0 22632 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0398_
timestamp 1667941163
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0399_
timestamp 1667941163
transform 1 0 12328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0400_
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0401_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0402_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0403_
timestamp 1667941163
transform 1 0 6716 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0404_
timestamp 1667941163
transform 1 0 12328 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0405_
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0406_
timestamp 1667941163
transform 1 0 12052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0407_
timestamp 1667941163
transform 1 0 6256 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0408_
timestamp 1667941163
transform 1 0 6900 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0409_
timestamp 1667941163
transform 1 0 4600 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0410_
timestamp 1667941163
transform 1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0411_
timestamp 1667941163
transform 1 0 11408 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 4416 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0414_
timestamp 1667941163
transform 1 0 4784 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0415_
timestamp 1667941163
transform 1 0 27600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0416_
timestamp 1667941163
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0417_
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 20608 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 28244 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0421_
timestamp 1667941163
transform 1 0 23828 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0423_
timestamp 1667941163
transform 1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 22908 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 24196 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0427_
timestamp 1667941163
transform 1 0 18124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0428_
timestamp 1667941163
transform 1 0 23276 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0429_
timestamp 1667941163
transform 1 0 23092 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0430_
timestamp 1667941163
transform 1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1667941163
transform 1 0 18032 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0434_
timestamp 1667941163
transform 1 0 27324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0435_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0436_
timestamp 1667941163
transform 1 0 27968 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 28520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 28612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0439_
timestamp 1667941163
transform 1 0 24104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 23276 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0441_
timestamp 1667941163
transform 1 0 23368 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 22448 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 25576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1667941163
transform 1 0 24104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0446_
timestamp 1667941163
transform 1 0 25484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0447_
timestamp 1667941163
transform 1 0 25944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448_
timestamp 1667941163
transform 1 0 22816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 19320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 23552 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 24196 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1667941163
transform 1 0 20792 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform 1 0 22172 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 22816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1667941163
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1667941163
transform 1 0 25024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 9936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0460_
timestamp 1667941163
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1667941163
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1667941163
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 23552 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 15456 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 16100 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 23184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 21712 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0473_
timestamp 1667941163
transform 1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 3220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 1840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform 1 0 17848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1667941163
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 7728 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 17204 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 12144 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 23736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 4968 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 18676 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 22448 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 9844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 15640 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 20424 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 22540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 18216 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 12420 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 6716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 10396 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 16008 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 18400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 23276 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 6532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 2668 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 6992 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 15088 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 14444 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 23092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 23092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 21804 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 17112 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 19780 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 3404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 18584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 2024 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 2852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 20608 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 9200 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 21528 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 23828 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 17848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 19872 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 14260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 15824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 19044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 16468 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 19596 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 23920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 23276 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 6532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 23276 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 20516 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 20516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 9292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 14904 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 9568 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 17112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 11776 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 11776 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 12880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 14076 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 18400 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 2300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 19596 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 4784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 25668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 12880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 27232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 8648 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 15364 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 26220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 5796 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 36708 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 9108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 31188 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 1840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 35880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 4968 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 23736 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 22448 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 21988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 22632 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 27140 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 35512 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 12328 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 28980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 21712 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 28612 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0653_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 29624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 29716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 4324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 9384 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 24748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 29900 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 5704 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 15088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 2668 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 25300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 22080 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 9016 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 32292 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 9384 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 6072 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0688_
timestamp 1667941163
transform 1 0 1840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 20700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 32292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 7360 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 31280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0696_
timestamp 1667941163
transform 1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 4048 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 15824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 5520 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 29256 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 5060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 28060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 28336 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 18400 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 25668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 23092 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 27784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 20240 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 29256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 27232 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 27784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 17940 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 26220 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 6624 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 31372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 3772 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 32016 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 4140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0727_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0728_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18032 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0729_
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 15824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 9936 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 16468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 6532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0740_
timestamp 1667941163
transform 1 0 13248 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 7176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 6440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 4232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0751_
timestamp 1667941163
transform 1 0 15824 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 6808 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 3956 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0762_
timestamp 1667941163
transform 1 0 14168 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0773_
timestamp 1667941163
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 24748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 10580 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0784_
timestamp 1667941163
transform 1 0 19596 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 4324 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 9292 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0795_
timestamp 1667941163
transform 1 0 13248 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 15916 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 23276 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 14904 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 9384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0806_
timestamp 1667941163
transform 1 0 18124 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 7268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 6624 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0817_
timestamp 1667941163
transform 1 0 12328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0828_
timestamp 1667941163
transform 1 0 18400 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 5428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 5612 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 5060 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 4784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 10488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0839_
timestamp 1667941163
transform 1 0 10672 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 9844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 10488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 10488 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 3128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 7820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 15640 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 10488 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 14720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0858_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 7360 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0862_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11224 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0863_
timestamp 1667941163
transform 1 0 7728 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0864_
timestamp 1667941163
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0865_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4508 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0866_
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 1656 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 4232 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0870_
timestamp 1667941163
transform 1 0 4048 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0871_
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0872_
timestamp 1667941163
transform 1 0 7912 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0873_
timestamp 1667941163
transform 1 0 11316 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0874_
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0875_
timestamp 1667941163
transform 1 0 5796 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 4232 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 3956 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0878_
timestamp 1667941163
transform 1 0 5428 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0879_
timestamp 1667941163
transform 1 0 3956 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0880_
timestamp 1667941163
transform 1 0 6532 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0881_
timestamp 1667941163
transform 1 0 4324 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0882_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1667941163
transform 1 0 9108 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 11224 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0885_
timestamp 1667941163
transform 1 0 6900 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0886_
timestamp 1667941163
transform 1 0 11684 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0887_
timestamp 1667941163
transform 1 0 9292 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0888_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0889_
timestamp 1667941163
transform 1 0 6808 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0890_
timestamp 1667941163
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1667941163
transform 1 0 13984 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0895_
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0896_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0897_
timestamp 1667941163
transform 1 0 11868 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0899_
timestamp 1667941163
transform 1 0 2392 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0902_
timestamp 1667941163
transform 1 0 6716 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0903_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0904_
timestamp 1667941163
transform 1 0 11868 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0905_
timestamp 1667941163
transform 1 0 10580 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 6624 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0907_
timestamp 1667941163
transform 1 0 4232 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 10304 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0910_
timestamp 1667941163
transform 1 0 11040 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0911_
timestamp 1667941163
transform 1 0 11960 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 1564 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0913_
timestamp 1667941163
transform 1 0 4140 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 1656 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0915_
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0916_
timestamp 1667941163
transform 1 0 7820 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform 1 0 8004 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 5888 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 4232 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 4232 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0921_
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0922_
timestamp 1667941163
transform 1 0 1564 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0923_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0924_
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 6808 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0927_
timestamp 1667941163
transform 1 0 11684 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0928_
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0929_
timestamp 1667941163
transform 1 0 11868 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 2024 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 4232 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1667941163
transform 1 0 14168 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0935_
timestamp 1667941163
transform 1 0 8280 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform 1 0 1656 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 2208 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 9384 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 11776 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0941_
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1667941163
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 5888 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 4140 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 3128 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0946_
timestamp 1667941163
transform 1 0 6164 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 4232 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 1656 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 4232 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 3956 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 5428 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 4232 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0954_
timestamp 1667941163
transform 1 0 11592 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0955_
timestamp 1667941163
transform 1 0 6532 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform 1 0 7176 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0957_
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0958_
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0959_
timestamp 1667941163
transform 1 0 7084 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1667941163
transform 1 0 9108 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0961_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0962_
timestamp 1667941163
transform 1 0 6624 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0963_
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0964_
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0965_
timestamp 1667941163
transform 1 0 7176 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0966_
timestamp 1667941163
transform 1 0 7820 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0967_
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0968_
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0969_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0970_
timestamp 1667941163
transform 1 0 1748 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0971_
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0972_
timestamp 1667941163
transform 1 0 13984 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0973_
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0974_
timestamp 1667941163
transform 1 0 11684 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0975_
timestamp 1667941163
transform 1 0 11684 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 35144 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1003_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 23552 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 32292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 30728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 32200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 33672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 25944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 4416 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 34224 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 27784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 32292 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 14168 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 32568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 7452 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 13156 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 18308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1024_
timestamp 1667941163
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 26036 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 35512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 30452 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1028_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1029_
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 5244 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 35328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 37812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1033_
timestamp 1667941163
transform 1 0 13156 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 35972 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1036_
timestamp 1667941163
transform 1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1037_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1042_
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1043_
timestamp 1667941163
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1044_
timestamp 1667941163
transform 1 0 18952 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1667941163
transform 1 0 36616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1046_
timestamp 1667941163
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1667941163
transform 1 0 35236 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1048_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1667941163
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1050_
timestamp 1667941163
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1667941163
transform 1 0 5704 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1052_
timestamp 1667941163
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1667941163
transform 1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1054_
timestamp 1667941163
transform 1 0 7176 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1056_
timestamp 1667941163
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 1667941163
transform 1 0 37812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1058_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12604 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 9936 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1060_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1060__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1061_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1062_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1063_
timestamp 1667941163
transform 1 0 14996 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1064_
timestamp 1667941163
transform 1 0 8004 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1065_
timestamp 1667941163
transform 1 0 21712 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1066_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1067_
timestamp 1667941163
transform 1 0 13984 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1068_
timestamp 1667941163
transform 1 0 24288 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1069_
timestamp 1667941163
transform 1 0 25208 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1070_
timestamp 1667941163
transform 1 0 14536 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1071_
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1072_
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1072__143
timestamp 1667941163
transform 1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1073_
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1074_
timestamp 1667941163
transform 1 0 10580 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1075_
timestamp 1667941163
transform 1 0 20056 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1076_
timestamp 1667941163
transform 1 0 1564 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1077_
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1078_
timestamp 1667941163
transform 1 0 15916 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1079_
timestamp 1667941163
transform 1 0 15364 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1080_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1081_
timestamp 1667941163
transform 1 0 16192 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1082_
timestamp 1667941163
transform 1 0 12420 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1083_
timestamp 1667941163
transform 1 0 18308 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1084_
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1084__144
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1085_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13892 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1086_
timestamp 1667941163
transform 1 0 13156 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1087_
timestamp 1667941163
transform 1 0 12420 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1088_
timestamp 1667941163
transform 1 0 8464 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1089_
timestamp 1667941163
transform 1 0 5796 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1090_
timestamp 1667941163
transform 1 0 13248 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1091_
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1092_
timestamp 1667941163
transform 1 0 12420 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1093_
timestamp 1667941163
transform 1 0 12420 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1094_
timestamp 1667941163
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1095_
timestamp 1667941163
transform 1 0 17204 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 19412 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1096__145
timestamp 1667941163
transform 1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1097_
timestamp 1667941163
transform 1 0 17296 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1098_
timestamp 1667941163
transform 1 0 18952 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1099_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1100_
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1101_
timestamp 1667941163
transform 1 0 19228 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 15548 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1103_
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1104_
timestamp 1667941163
transform 1 0 16836 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 14352 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1106_
timestamp 1667941163
transform 1 0 16560 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1107_
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1108_
timestamp 1667941163
transform 1 0 19228 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1108__146
timestamp 1667941163
transform 1 0 18584 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1109_
timestamp 1667941163
transform 1 0 16928 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1110_
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1112_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1113_
timestamp 1667941163
transform 1 0 17296 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1114_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1115_
timestamp 1667941163
transform 1 0 16928 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1116_
timestamp 1667941163
transform 1 0 18124 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 18400 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1118_
timestamp 1667941163
transform 1 0 9200 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 1748 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1120__147
timestamp 1667941163
transform 1 0 2760 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1120_
timestamp 1667941163
transform 1 0 2116 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1121_
timestamp 1667941163
transform 1 0 20332 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1122_
timestamp 1667941163
transform 1 0 13984 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1123_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1124_
timestamp 1667941163
transform 1 0 7084 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1125_
timestamp 1667941163
transform 1 0 18492 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1126_
timestamp 1667941163
transform 1 0 1656 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1127_
timestamp 1667941163
transform 1 0 4416 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1128_
timestamp 1667941163
transform 1 0 20056 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1129_
timestamp 1667941163
transform 1 0 18308 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1130_
timestamp 1667941163
transform 1 0 15088 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1132_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1133__148
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1133_
timestamp 1667941163
transform 1 0 19228 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 19596 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1136_
timestamp 1667941163
transform 1 0 19596 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 20240 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 17664 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 19412 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1140_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 17112 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1142_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1143_
timestamp 1667941163
transform 1 0 7452 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 17112 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1145__149
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1145_
timestamp 1667941163
transform 1 0 13616 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform 1 0 18492 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 17388 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 21344 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1150_
timestamp 1667941163
transform 1 0 2300 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1151_
timestamp 1667941163
transform 1 0 8648 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1152_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 6532 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1154_
timestamp 1667941163
transform 1 0 13892 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1155_
timestamp 1667941163
transform 1 0 17940 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 18032 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1157__150
timestamp 1667941163
transform 1 0 24104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1157_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1158_
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1159_
timestamp 1667941163
transform 1 0 14260 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 13616 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 15272 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1162_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 1656 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1166_
timestamp 1667941163
transform 1 0 10028 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1167_
timestamp 1667941163
transform 1 0 11960 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 11224 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1169__151
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1169_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 9936 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform 1 0 24748 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1173_
timestamp 1667941163
transform 1 0 19688 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1174_
timestamp 1667941163
transform 1 0 14076 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1175_
timestamp 1667941163
transform 1 0 17020 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 9936 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1177_
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1178_
timestamp 1667941163
transform 1 0 16100 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1179_
timestamp 1667941163
transform 1 0 16468 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1180__152
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1180_
timestamp 1667941163
transform 1 0 10396 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 20516 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 17664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1184_
timestamp 1667941163
transform 1 0 13984 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1185_
timestamp 1667941163
transform 1 0 14628 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1186_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1187_
timestamp 1667941163
transform 1 0 16560 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1188_
timestamp 1667941163
transform 1 0 4968 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1188__153
timestamp 1667941163
transform 1 0 4140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1189_
timestamp 1667941163
transform 1 0 19872 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 16560 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 16836 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1192_
timestamp 1667941163
transform 1 0 17204 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1193_
timestamp 1667941163
transform 1 0 17940 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1194_
timestamp 1667941163
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1195_
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1196__154
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1197_
timestamp 1667941163
transform 1 0 7360 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1198_
timestamp 1667941163
transform 1 0 15548 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1200_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1201_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 4600 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1203__155
timestamp 1667941163
transform 1 0 6808 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1203_
timestamp 1667941163
transform 1 0 6624 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1204_
timestamp 1667941163
transform 1 0 4324 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1205_
timestamp 1667941163
transform 1 0 11040 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1206_
timestamp 1667941163
transform 1 0 7912 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1207_
timestamp 1667941163
transform 1 0 9844 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1209__156
timestamp 1667941163
transform 1 0 25944 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 24932 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 14352 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1211_
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 20424 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 23092 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 19688 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1215__157
timestamp 1667941163
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 16468 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1217_
timestamp 1667941163
transform 1 0 15548 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1667941163
transform 1 0 21160 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1219_
timestamp 1667941163
transform 1 0 21252 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform 1 0 21344 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1221__158
timestamp 1667941163
transform 1 0 20700 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1222_
timestamp 1667941163
transform 1 0 18032 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1223_
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1224_
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1225_
timestamp 1667941163
transform 1 0 19044 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1226_
timestamp 1667941163
transform 1 0 24472 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1227__159
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1667941163
transform 1 0 25760 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1228_
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1667941163
transform 1 0 23000 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1230_
timestamp 1667941163
transform 1 0 22356 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1667941163
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1232_
timestamp 1667941163
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1233_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1233__160
timestamp 1667941163
transform 1 0 26680 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1234_
timestamp 1667941163
transform 1 0 20792 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1235_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1236_
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1237_
timestamp 1667941163
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1238_
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1239__161
timestamp 1667941163
transform 1 0 21712 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1239_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1240_
timestamp 1667941163
transform 1 0 21804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1241_
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1242_
timestamp 1667941163
transform 1 0 16928 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1243_
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1244__162
timestamp 1667941163
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1244_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1245_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1246_
timestamp 1667941163
transform 1 0 26128 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1247_
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1248__163
timestamp 1667941163
transform 1 0 3128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1248_
timestamp 1667941163
transform 1 0 3220 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1249_
timestamp 1667941163
transform 1 0 9844 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1250_
timestamp 1667941163
transform 1 0 3128 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1251_
timestamp 1667941163
transform 1 0 7820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1252_
timestamp 1667941163
transform 1 0 9108 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1252__164
timestamp 1667941163
transform 1 0 8004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1253_
timestamp 1667941163
transform 1 0 10948 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1254_
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1255_
timestamp 1667941163
transform 1 0 12420 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1256__165
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1256_
timestamp 1667941163
transform 1 0 23092 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1257_
timestamp 1667941163
transform 1 0 11960 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1258_
timestamp 1667941163
transform 1 0 21068 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1259_
timestamp 1667941163
transform 1 0 12696 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1260_
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1260__166
timestamp 1667941163
transform 1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1261_
timestamp 1667941163
transform 1 0 10672 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1262_
timestamp 1667941163
transform 1 0 25852 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1263_
timestamp 1667941163
transform 1 0 3128 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4232 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 6532 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 9660 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 13892 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 9936 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 14352 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 3956 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 3956 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 7636 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 14168 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 10028 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 5796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 1564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 38088 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 3956 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 12972 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 38088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 35328 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 37444 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 38088 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 38088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 15548 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 33028 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 25208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1667941163
transform 1 0 30912 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 25024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 6532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 6716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1667941163
transform 1 0 2852 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1667941163
transform 1 0 3128 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1667941163
transform 1 0 37260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 14260 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1667941163
transform 1 0 2116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1667941163
transform 1 0 37444 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1667941163
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1667941163
transform 1 0 37444 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 38088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 2300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1667941163
transform 1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 2852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 38088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 37996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 17480 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 9108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 21988 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  sb_4__1__141
timestamp 1667941163
transform 1 0 25852 0 -1 4352
box -38 -48 314 592
<< labels >>
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 2 nsew signal input
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 3 nsew signal input
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 4 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 5 nsew signal input
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 6 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 8 nsew signal input
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 9 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 ccff_head
port 10 nsew signal input
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 12 nsew signal input
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 13 nsew signal input
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 14 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 15 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 16 nsew signal input
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 17 nsew signal input
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 18 nsew signal input
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 19 nsew signal input
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_left_in[17]
port 20 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 21 nsew signal input
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 22 nsew signal input
flabel metal3 s 39200 27888 39800 28008 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 23 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 24 nsew signal input
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 25 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 26 nsew signal input
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 27 nsew signal input
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 28 nsew signal input
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 29 nsew signal input
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 chanx_left_in[9]
port 30 nsew signal input
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 31 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 32 nsew signal tristate
flabel metal3 s 39200 12928 39800 13048 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 33 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 34 nsew signal tristate
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 35 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 36 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 37 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 38 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 39 nsew signal tristate
flabel metal3 s 39200 16328 39800 16448 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 40 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 41 nsew signal tristate
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 42 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 43 nsew signal tristate
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 44 nsew signal tristate
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 45 nsew signal tristate
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 46 nsew signal tristate
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 47 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 48 nsew signal tristate
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 49 nsew signal tristate
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 17406 39200 17462 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal2 s 14186 39200 14242 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 98 nsew signal input
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_top_in[2]
port 99 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_top_in[3]
port 100 nsew signal input
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_top_in[4]
port 101 nsew signal input
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_top_in[5]
port 102 nsew signal input
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 103 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_in[7]
port 104 nsew signal input
flabel metal3 s 39200 9528 39800 9648 0 FreeSans 480 0 0 0 chany_top_in[8]
port 105 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_in[9]
port 106 nsew signal input
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_top_out[0]
port 107 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_out[10]
port 108 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 109 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_top_out[12]
port 110 nsew signal tristate
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_top_out[13]
port 111 nsew signal tristate
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chany_top_out[14]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_top_out[15]
port 113 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 114 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 115 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chany_top_out[18]
port 116 nsew signal tristate
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 117 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 126 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 127 nsew signal input
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 128 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 129 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 pReset
port 130 nsew signal input
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 prog_clk
port 131 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 132 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 133 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 137 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 138 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 139 nsew signal input
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 140 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 141 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 11500 10778 11500 10778 0 _0000_
rlabel metal1 14904 15334 14904 15334 0 _0001_
rlabel metal1 7774 4998 7774 4998 0 _0002_
rlabel metal1 5842 8398 5842 8398 0 _0003_
rlabel metal1 6762 4658 6762 4658 0 _0004_
rlabel metal1 5520 7310 5520 7310 0 _0005_
rlabel via2 5382 12189 5382 12189 0 _0006_
rlabel metal2 10718 9588 10718 9588 0 _0007_
rlabel metal2 1794 10880 1794 10880 0 _0008_
rlabel metal2 12834 6562 12834 6562 0 _0009_
rlabel metal1 5244 7854 5244 7854 0 _0010_
rlabel metal1 6302 3094 6302 3094 0 _0011_
rlabel metal1 7268 2822 7268 2822 0 _0012_
rlabel metal2 13110 6086 13110 6086 0 _0013_
rlabel metal1 4830 3944 4830 3944 0 _0014_
rlabel metal2 25530 3757 25530 3757 0 _0015_
rlabel metal1 10810 2278 10810 2278 0 _0016_
rlabel metal2 15502 2142 15502 2142 0 _0017_
rlabel metal1 6079 18734 6079 18734 0 _0018_
rlabel metal1 3503 17578 3503 17578 0 _0019_
rlabel via2 9522 14331 9522 14331 0 _0020_
rlabel metal1 8043 13974 8043 13974 0 _0021_
rlabel metal2 7866 14824 7866 14824 0 _0022_
rlabel metal2 10442 4488 10442 4488 0 _0023_
rlabel metal2 12282 4403 12282 4403 0 _0024_
rlabel metal1 9706 8534 9706 8534 0 _0025_
rlabel metal1 15962 16762 15962 16762 0 _0026_
rlabel metal1 8464 7718 8464 7718 0 _0027_
rlabel metal1 13432 3706 13432 3706 0 _0028_
rlabel via2 4094 12869 4094 12869 0 _0029_
rlabel metal1 15088 8602 15088 8602 0 _0030_
rlabel metal1 14444 16014 14444 16014 0 _0031_
rlabel metal2 11270 13022 11270 13022 0 _0032_
rlabel metal1 9614 11560 9614 11560 0 _0033_
rlabel metal1 13570 4794 13570 4794 0 _0034_
rlabel metal2 23414 3213 23414 3213 0 _0035_
rlabel metal1 3588 3366 3588 3366 0 _0036_
rlabel metal2 17618 5287 17618 5287 0 _0037_
rlabel metal1 15739 4590 15739 4590 0 _0038_
rlabel metal2 22034 4352 22034 4352 0 _0039_
rlabel via2 22770 4267 22770 4267 0 _0040_
rlabel metal1 6302 11662 6302 11662 0 _0041_
rlabel metal1 6624 4794 6624 4794 0 _0042_
rlabel metal1 20010 1904 20010 1904 0 _0043_
rlabel metal2 17986 2176 17986 2176 0 _0044_
rlabel metal2 7222 2992 7222 2992 0 _0045_
rlabel metal1 5382 3162 5382 3162 0 _0046_
rlabel metal2 5290 8704 5290 8704 0 _0047_
rlabel metal1 7827 7786 7827 7786 0 _0048_
rlabel metal1 5106 3094 5106 3094 0 _0049_
rlabel metal1 6992 2958 6992 2958 0 _0050_
rlabel via2 16054 3179 16054 3179 0 _0051_
rlabel metal1 16974 3502 16974 3502 0 _0052_
rlabel metal1 3503 16558 3503 16558 0 _0053_
rlabel metal1 5704 23494 5704 23494 0 _0054_
rlabel metal3 5727 21284 5727 21284 0 _0055_
rlabel metal1 5244 24582 5244 24582 0 _0056_
rlabel metal2 5612 17068 5612 17068 0 _0057_
rlabel metal1 9706 14246 9706 14246 0 _0058_
rlabel metal1 13432 16762 13432 16762 0 _0059_
rlabel metal1 7031 18326 7031 18326 0 _0060_
rlabel metal1 7912 3638 7912 3638 0 _0061_
rlabel via2 9614 9605 9614 9605 0 _0062_
rlabel metal1 12183 14314 12183 14314 0 _0063_
rlabel metal2 15594 15657 15594 15657 0 _0064_
rlabel metal2 9890 6766 9890 6766 0 _0065_
rlabel metal1 15410 14042 15410 14042 0 _0066_
rlabel metal2 15410 3655 15410 3655 0 _0067_
rlabel metal2 8510 6120 8510 6120 0 _0068_
rlabel metal2 11086 14688 11086 14688 0 _0069_
rlabel metal1 6716 9146 6716 9146 0 _0070_
rlabel metal2 10626 8262 10626 8262 0 _0071_
rlabel metal2 21666 6392 21666 6392 0 _0072_
rlabel metal2 3220 15572 3220 15572 0 _0073_
rlabel metal1 10994 15096 10994 15096 0 _0074_
rlabel via3 3381 17884 3381 17884 0 _0075_
rlabel metal1 4002 18394 4002 18394 0 _0076_
rlabel metal1 15916 2822 15916 2822 0 _0077_
rlabel metal1 15318 16150 15318 16150 0 _0078_
rlabel metal1 10718 16218 10718 16218 0 _0079_
rlabel metal1 14352 10438 14352 10438 0 _0080_
rlabel metal1 4370 14790 4370 14790 0 _0081_
rlabel metal1 3503 15402 3503 15402 0 _0082_
rlabel metal1 15548 13158 15548 13158 0 _0083_
rlabel metal2 10074 18462 10074 18462 0 _0084_
rlabel metal1 9016 10778 9016 10778 0 _0085_
rlabel metal1 9154 17129 9154 17129 0 _0086_
rlabel metal1 7038 13974 7038 13974 0 _0087_
rlabel metal1 7452 2618 7452 2618 0 _0088_
rlabel metal3 13892 1564 13892 1564 0 _0089_
rlabel metal1 8464 3162 8464 3162 0 _0090_
rlabel metal1 10350 2618 10350 2618 0 _0091_
rlabel metal3 9108 12512 9108 12512 0 _0092_
rlabel metal2 5106 19618 5106 19618 0 _0093_
rlabel metal1 4423 14314 4423 14314 0 _0094_
rlabel metal1 8595 11798 8595 11798 0 _0095_
rlabel metal1 8280 3366 8280 3366 0 _0096_
rlabel metal1 8464 13226 8464 13226 0 _0097_
rlabel metal2 7222 13498 7222 13498 0 _0098_
rlabel metal1 5803 16150 5803 16150 0 _0099_
rlabel metal1 4416 21930 4416 21930 0 _0100_
rlabel via1 6762 14331 6762 14331 0 _0101_
rlabel metal2 5014 16201 5014 16201 0 _0102_
rlabel via2 7843 21828 7843 21828 0 _0103_
rlabel metal1 8556 6630 8556 6630 0 _0104_
rlabel metal2 15226 8568 15226 8568 0 _0105_
rlabel metal3 20148 7480 20148 7480 0 _0106_
rlabel metal1 4830 2958 4830 2958 0 _0107_
rlabel metal2 19274 2176 19274 2176 0 _0108_
rlabel metal2 20470 4624 20470 4624 0 _0109_
rlabel metal1 19090 2074 19090 2074 0 _0110_
rlabel metal2 15042 4743 15042 4743 0 _0111_
rlabel metal1 7222 3162 7222 3162 0 _0112_
rlabel metal2 18538 15504 18538 15504 0 _0113_
rlabel metal2 12466 13197 12466 13197 0 _0114_
rlabel metal2 13754 10744 13754 10744 0 _0115_
rlabel metal2 14674 7820 14674 7820 0 _0116_
rlabel metal2 11546 9027 11546 9027 0 _0117_
rlabel metal1 9384 2550 9384 2550 0 _0118_
rlabel metal2 16146 6460 16146 6460 0 _0119_
rlabel metal1 14168 7446 14168 7446 0 _0120_
rlabel metal1 1702 10608 1702 10608 0 _0121_
rlabel metal1 8418 2380 8418 2380 0 _0122_
rlabel metal2 21114 13175 21114 13175 0 _0123_
rlabel metal1 19274 7854 19274 7854 0 _0124_
rlabel metal1 7498 3026 7498 3026 0 _0125_
rlabel metal2 9062 9503 9062 9503 0 _0126_
rlabel metal1 15594 13940 15594 13940 0 _0127_
rlabel metal1 10764 23698 10764 23698 0 _0128_
rlabel metal1 26404 19822 26404 19822 0 _0129_
rlabel metal2 12466 22474 12466 22474 0 _0130_
rlabel metal2 24794 10506 24794 10506 0 _0131_
rlabel metal2 12282 26826 12282 26826 0 _0132_
rlabel metal1 7130 26384 7130 26384 0 _0133_
rlabel metal2 11086 27132 11086 27132 0 _0134_
rlabel metal2 5014 24378 5014 24378 0 _0135_
rlabel metal2 20838 16388 20838 16388 0 _0136_
rlabel metal1 29118 16116 29118 16116 0 _0137_
rlabel metal1 23368 15470 23368 15470 0 _0138_
rlabel metal1 24150 18394 24150 18394 0 _0139_
rlabel metal2 23322 23290 23322 23290 0 _0140_
rlabel metal1 21758 19346 21758 19346 0 _0141_
rlabel metal2 27370 14076 27370 14076 0 _0142_
rlabel metal2 28842 15164 28842 15164 0 _0143_
rlabel metal1 23046 13294 23046 13294 0 _0144_
rlabel metal2 24610 9350 24610 9350 0 _0145_
rlabel metal2 26174 11322 26174 11322 0 _0146_
rlabel metal1 19504 25874 19504 25874 0 _0147_
rlabel metal1 24150 24786 24150 24786 0 _0148_
rlabel metal1 23046 26316 23046 26316 0 _0149_
rlabel metal2 13340 8602 13340 8602 0 _0150_
rlabel metal2 20378 4420 20378 4420 0 _0151_
rlabel metal2 26450 6086 26450 6086 0 _0152_
rlabel metal1 16330 20876 16330 20876 0 _0153_
rlabel metal2 23414 18700 23414 18700 0 _0154_
rlabel metal2 25070 18564 25070 18564 0 _0155_
rlabel metal1 18262 11118 18262 11118 0 _0156_
rlabel metal1 16008 2414 16008 2414 0 _0157_
rlabel metal1 7498 2414 7498 2414 0 _0158_
rlabel metal2 12926 15266 12926 15266 0 _0159_
rlabel metal1 9936 20774 9936 20774 0 _0160_
rlabel metal2 17066 15198 17066 15198 0 _0161_
rlabel metal2 9338 22440 9338 22440 0 _0162_
rlabel metal1 25576 16218 25576 16218 0 _0163_
rlabel metal1 15364 22406 15364 22406 0 _0164_
rlabel metal1 8510 20502 8510 20502 0 _0165_
rlabel via2 21942 11067 21942 11067 0 _0166_
rlabel metal2 14490 20298 14490 20298 0 _0167_
rlabel metal1 14214 15096 14214 15096 0 _0168_
rlabel metal1 25162 17238 25162 17238 0 _0169_
rlabel metal1 25346 21658 25346 21658 0 _0170_
rlabel metal1 13478 8908 13478 8908 0 _0171_
rlabel metal1 19458 3162 19458 3162 0 _0172_
rlabel metal1 14582 6834 14582 6834 0 _0173_
rlabel metal2 21298 12274 21298 12274 0 _0174_
rlabel metal1 5980 14586 5980 14586 0 _0175_
rlabel metal1 20286 11016 20286 11016 0 _0176_
rlabel metal1 2254 24854 2254 24854 0 _0177_
rlabel metal1 1978 19414 1978 19414 0 _0178_
rlabel metal1 16284 26282 16284 26282 0 _0179_
rlabel metal1 13662 14280 13662 14280 0 _0180_
rlabel metal1 22172 15130 22172 15130 0 _0181_
rlabel metal1 17848 21590 17848 21590 0 _0182_
rlabel metal1 12650 20808 12650 20808 0 _0183_
rlabel metal2 17250 19720 17250 19720 0 _0184_
rlabel metal1 16054 19482 16054 19482 0 _0185_
rlabel metal2 14122 25262 14122 25262 0 _0186_
rlabel metal1 13938 21590 13938 21590 0 _0187_
rlabel metal2 12650 25704 12650 25704 0 _0188_
rlabel metal1 8694 23800 8694 23800 0 _0189_
rlabel metal1 5980 22610 5980 22610 0 _0190_
rlabel metal1 13938 27030 13938 27030 0 _0191_
rlabel metal1 14306 26248 14306 26248 0 _0192_
rlabel metal2 12650 23086 12650 23086 0 _0193_
rlabel metal1 12650 23800 12650 23800 0 _0194_
rlabel metal2 20654 6324 20654 6324 0 _0195_
rlabel metal2 16422 10098 16422 10098 0 _0196_
rlabel metal1 22126 8058 22126 8058 0 _0197_
rlabel metal1 20470 5752 20470 5752 0 _0198_
rlabel metal2 20654 16456 20654 16456 0 _0199_
rlabel metal1 11408 20502 11408 20502 0 _0200_
rlabel metal2 21666 7650 21666 7650 0 _0201_
rlabel metal1 21114 5746 21114 5746 0 _0202_
rlabel metal1 21942 6120 21942 6120 0 _0203_
rlabel metal1 20095 3128 20095 3128 0 _0204_
rlabel metal1 16974 5032 16974 5032 0 _0205_
rlabel metal2 14582 3570 14582 3570 0 _0206_
rlabel metal1 15732 14586 15732 14586 0 _0207_
rlabel metal1 16284 17850 16284 17850 0 _0208_
rlabel metal1 19458 16184 19458 16184 0 _0209_
rlabel metal1 19596 18938 19596 18938 0 _0210_
rlabel metal1 14490 18632 14490 18632 0 _0211_
rlabel metal1 15410 23018 15410 23018 0 _0212_
rlabel metal1 19826 15402 19826 15402 0 _0213_
rlabel metal1 17710 14314 17710 14314 0 _0214_
rlabel metal2 21758 11424 21758 11424 0 _0215_
rlabel metal1 21114 13498 21114 13498 0 _0216_
rlabel metal2 19182 21760 19182 21760 0 _0217_
rlabel metal1 21712 7446 21712 7446 0 _0218_
rlabel metal2 9430 21080 9430 21080 0 _0219_
rlabel metal1 1978 22712 1978 22712 0 _0220_
rlabel metal1 2254 26282 2254 26282 0 _0221_
rlabel metal1 20424 12614 20424 12614 0 _0222_
rlabel via2 9338 16779 9338 16779 0 _0223_
rlabel metal2 20746 10472 20746 10472 0 _0224_
rlabel metal1 7360 21590 7360 21590 0 _0225_
rlabel metal2 18722 13022 18722 13022 0 _0226_
rlabel metal2 1886 23630 1886 23630 0 _0227_
rlabel metal1 4692 21590 4692 21590 0 _0228_
rlabel metal1 20562 10710 20562 10710 0 _0229_
rlabel metal2 18906 10676 18906 10676 0 _0230_
rlabel metal1 9844 3706 9844 3706 0 _0231_
rlabel metal1 18814 3162 18814 3162 0 _0232_
rlabel metal1 19918 4658 19918 4658 0 _0233_
rlabel metal1 20332 4046 20332 4046 0 _0234_
rlabel metal1 20010 13498 20010 13498 0 _0235_
rlabel metal1 16514 17238 16514 17238 0 _0236_
rlabel metal1 20102 5270 20102 5270 0 _0237_
rlabel metal1 20470 7752 20470 7752 0 _0238_
rlabel metal1 17894 3400 17894 3400 0 _0239_
rlabel metal1 19642 5644 19642 5644 0 _0240_
rlabel metal2 17342 15810 17342 15810 0 _0241_
rlabel metal1 18354 5304 18354 5304 0 _0242_
rlabel metal1 15732 17306 15732 17306 0 _0243_
rlabel metal2 7682 20876 7682 20876 0 _0244_
rlabel metal2 18170 20400 18170 20400 0 _0245_
rlabel metal2 13846 22916 13846 22916 0 _0246_
rlabel metal2 18722 14110 18722 14110 0 _0247_
rlabel metal2 17618 23902 17618 23902 0 _0248_
rlabel metal1 21574 19720 21574 19720 0 _0249_
rlabel metal1 10948 20570 10948 20570 0 _0250_
rlabel metal2 2530 15266 2530 15266 0 _0251_
rlabel metal1 9338 21590 9338 21590 0 _0252_
rlabel metal1 14904 27098 14904 27098 0 _0253_
rlabel metal1 6946 20502 6946 20502 0 _0254_
rlabel metal1 9522 12886 9522 12886 0 _0255_
rlabel metal1 18354 4794 18354 4794 0 _0256_
rlabel metal1 20194 8024 20194 8024 0 _0257_
rlabel metal1 19734 9962 19734 9962 0 _0258_
rlabel metal2 2622 24854 2622 24854 0 _0259_
rlabel metal1 14536 20842 14536 20842 0 _0260_
rlabel metal1 14950 23766 14950 23766 0 _0261_
rlabel metal2 15502 20910 15502 20910 0 _0262_
rlabel metal2 13478 12937 13478 12937 0 _0263_
rlabel metal1 14950 3162 14950 3162 0 _0264_
rlabel metal1 1610 23052 1610 23052 0 _0265_
rlabel metal1 15134 22678 15134 22678 0 _0266_
rlabel metal1 10258 19448 10258 19448 0 _0267_
rlabel metal2 12190 20536 12190 20536 0 _0268_
rlabel metal2 11454 25432 11454 25432 0 _0269_
rlabel metal1 16928 24854 16928 24854 0 _0270_
rlabel metal2 10166 23902 10166 23902 0 _0271_
rlabel metal2 24978 19550 24978 19550 0 _0272_
rlabel metal1 19642 22984 19642 22984 0 _0273_
rlabel metal1 19964 21590 19964 21590 0 _0274_
rlabel metal1 15042 19414 15042 19414 0 _0275_
rlabel metal1 17250 25160 17250 25160 0 _0276_
rlabel metal1 10212 24106 10212 24106 0 _0277_
rlabel metal2 20562 21522 20562 21522 0 _0278_
rlabel metal1 16514 10030 16514 10030 0 _0279_
rlabel metal1 11270 11288 11270 11288 0 _0280_
rlabel metal1 10074 16558 10074 16558 0 _0281_
rlabel metal1 21298 6800 21298 6800 0 _0282_
rlabel metal1 20286 2278 20286 2278 0 _0283_
rlabel metal1 13708 11254 13708 11254 0 _0284_
rlabel metal1 13294 6120 13294 6120 0 _0285_
rlabel metal1 17572 2618 17572 2618 0 _0286_
rlabel metal2 20930 8704 20930 8704 0 _0287_
rlabel metal2 17894 8194 17894 8194 0 _0288_
rlabel metal1 5152 23494 5152 23494 0 _0289_
rlabel metal1 20608 8534 20608 8534 0 _0290_
rlabel metal2 21298 4828 21298 4828 0 _0291_
rlabel metal2 18814 7684 18814 7684 0 _0292_
rlabel metal2 18446 5304 18446 5304 0 _0293_
rlabel via2 19366 8789 19366 8789 0 _0294_
rlabel metal1 15732 18258 15732 18258 0 _0295_
rlabel metal2 9982 11407 9982 11407 0 _0296_
rlabel metal1 19090 11832 19090 11832 0 _0297_
rlabel metal2 7590 21352 7590 21352 0 _0298_
rlabel metal2 17710 3621 17710 3621 0 _0299_
rlabel metal1 17204 10642 17204 10642 0 _0300_
rlabel metal2 20378 12954 20378 12954 0 _0301_
rlabel metal1 17526 11798 17526 11798 0 _0302_
rlabel metal2 4830 21488 4830 21488 0 _0303_
rlabel metal1 4968 23290 4968 23290 0 _0304_
rlabel metal1 5014 20536 5014 20536 0 _0305_
rlabel metal1 5290 21862 5290 21862 0 _0306_
rlabel metal1 6210 22746 6210 22746 0 _0307_
rlabel metal1 10948 22746 10948 22746 0 _0308_
rlabel metal2 23230 18530 23230 18530 0 _0309_
rlabel metal1 25162 18836 25162 18836 0 _0310_
rlabel metal2 16146 21284 16146 21284 0 _0311_
rlabel metal2 23966 19584 23966 19584 0 _0312_
rlabel metal1 20792 13362 20792 13362 0 _0313_
rlabel metal2 23690 21012 23690 21012 0 _0314_
rlabel metal2 20562 5576 20562 5576 0 _0315_
rlabel metal1 25392 6426 25392 6426 0 _0316_
rlabel metal1 13708 13226 13708 13226 0 _0317_
rlabel metal1 20976 4794 20976 4794 0 _0318_
rlabel metal1 22126 6868 22126 6868 0 _0319_
rlabel metal2 21482 8704 21482 8704 0 _0320_
rlabel metal2 22218 24718 22218 24718 0 _0321_
rlabel metal2 22862 25772 22862 25772 0 _0322_
rlabel metal1 18814 24786 18814 24786 0 _0323_
rlabel metal1 20470 24072 20470 24072 0 _0324_
rlabel metal2 20194 25534 20194 25534 0 _0325_
rlabel metal2 19274 23868 19274 23868 0 _0326_
rlabel metal1 24702 9452 24702 9452 0 _0327_
rlabel metal2 25990 10812 25990 10812 0 _0328_
rlabel metal2 22494 13668 22494 13668 0 _0329_
rlabel metal1 23736 8398 23736 8398 0 _0330_
rlabel metal2 22586 11084 22586 11084 0 _0331_
rlabel metal1 22218 9486 22218 9486 0 _0332_
rlabel metal1 26680 13906 26680 13906 0 _0333_
rlabel metal1 27370 14892 27370 14892 0 _0334_
rlabel metal1 21160 17714 21160 17714 0 _0335_
rlabel metal2 24794 14620 24794 14620 0 _0336_
rlabel metal1 26358 13328 26358 13328 0 _0337_
rlabel metal2 18354 17340 18354 17340 0 _0338_
rlabel metal1 24058 20570 24058 20570 0 _0339_
rlabel metal1 22678 22950 22678 22950 0 _0340_
rlabel metal1 22080 15470 22080 15470 0 _0341_
rlabel metal2 23966 16898 23966 16898 0 _0342_
rlabel metal1 17572 20434 17572 20434 0 _0343_
rlabel metal1 20424 13838 20424 13838 0 _0344_
rlabel metal2 24794 15708 24794 15708 0 _0345_
rlabel metal1 19964 14450 19964 14450 0 _0346_
rlabel metal2 27738 16422 27738 16422 0 _0347_
rlabel metal1 19826 14994 19826 14994 0 _0348_
rlabel metal1 4462 21862 4462 21862 0 _0349_
rlabel metal2 10074 26588 10074 26588 0 _0350_
rlabel metal1 4002 23766 4002 23766 0 _0351_
rlabel metal2 8050 26316 8050 26316 0 _0352_
rlabel metal2 9338 25670 9338 25670 0 _0353_
rlabel metal2 11178 26282 11178 26282 0 _0354_
rlabel metal1 7820 27030 7820 27030 0 _0355_
rlabel metal1 12604 25330 12604 25330 0 _0356_
rlabel metal1 23414 9962 23414 9962 0 _0357_
rlabel metal2 12282 21726 12282 21726 0 _0358_
rlabel metal1 21298 9928 21298 9928 0 _0359_
rlabel metal1 12558 19414 12558 19414 0 _0360_
rlabel metal2 25806 20264 25806 20264 0 _0361_
rlabel metal1 10626 23494 10626 23494 0 _0362_
rlabel metal2 26266 21352 26266 21352 0 _0363_
rlabel metal1 3358 20536 3358 20536 0 _0364_
rlabel metal3 1234 28628 1234 28628 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 5934 37230 5934 37230 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 12926 2506 12926 2506 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 19366 1860 19366 1860 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1050 26588 1050 26588 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 11086 6953 11086 6953 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel via2 38318 30685 38318 30685 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 11730 493 11730 493 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 25346 37230 25346 37230 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 38318 8347 38318 8347 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal3 1050 748 1050 748 0 ccff_head
rlabel via2 38226 35445 38226 35445 0 ccff_tail
rlabel metal3 1717 19108 1717 19108 0 chanx_left_in[0]
rlabel metal1 26910 37230 26910 37230 0 chanx_left_in[10]
rlabel via2 3542 23205 3542 23205 0 chanx_left_in[11]
rlabel metal1 12834 37230 12834 37230 0 chanx_left_in[12]
rlabel metal2 38318 11033 38318 11033 0 chanx_left_in[13]
rlabel metal2 28382 1588 28382 1588 0 chanx_left_in[14]
rlabel metal1 4738 37230 4738 37230 0 chanx_left_in[15]
rlabel metal2 36110 38022 36110 38022 0 chanx_left_in[16]
rlabel metal1 37536 35054 37536 35054 0 chanx_left_in[17]
rlabel metal3 751 5508 751 5508 0 chanx_left_in[18]
rlabel metal2 20654 1588 20654 1588 0 chanx_left_in[1]
rlabel metal2 38318 27999 38318 27999 0 chanx_left_in[2]
rlabel metal2 38318 12563 38318 12563 0 chanx_left_in[3]
rlabel metal1 15640 37230 15640 37230 0 chanx_left_in[4]
rlabel metal2 39330 1860 39330 1860 0 chanx_left_in[5]
rlabel metal1 33074 37230 33074 37230 0 chanx_left_in[6]
rlabel metal2 17434 1214 17434 1214 0 chanx_left_in[7]
rlabel metal1 3726 37230 3726 37230 0 chanx_left_in[8]
rlabel metal2 10902 527 10902 527 0 chanx_left_in[9]
rlabel metal2 2806 14875 2806 14875 0 chanx_left_out[0]
rlabel metal2 25162 1520 25162 1520 0 chanx_left_out[10]
rlabel metal2 38226 13073 38226 13073 0 chanx_left_out[11]
rlabel via2 38226 27285 38226 27285 0 chanx_left_out[12]
rlabel metal2 34822 1520 34822 1520 0 chanx_left_out[13]
rlabel metal1 32384 37094 32384 37094 0 chanx_left_out[15]
rlabel metal1 20148 37094 20148 37094 0 chanx_left_out[16]
rlabel metal2 33534 1520 33534 1520 0 chanx_left_out[17]
rlabel via2 38226 16405 38226 16405 0 chanx_left_out[18]
rlabel metal1 7912 37094 7912 37094 0 chanx_left_out[1]
rlabel metal2 38226 23953 38226 23953 0 chanx_left_out[2]
rlabel metal1 16928 36890 16928 36890 0 chanx_left_out[3]
rlabel via2 38226 32725 38226 32725 0 chanx_left_out[4]
rlabel metal3 1234 4148 1234 4148 0 chanx_left_out[5]
rlabel metal2 38226 17901 38226 17901 0 chanx_left_out[6]
rlabel metal3 1234 31348 1234 31348 0 chanx_left_out[7]
rlabel metal3 1234 35428 1234 35428 0 chanx_left_out[8]
rlabel metal2 38226 32113 38226 32113 0 chanx_left_out[9]
rlabel metal1 37674 4182 37674 4182 0 chany_bottom_in[0]
rlabel metal1 21666 37298 21666 37298 0 chany_bottom_in[10]
rlabel metal1 19550 37230 19550 37230 0 chany_bottom_in[11]
rlabel metal2 30958 38260 30958 38260 0 chany_bottom_in[12]
rlabel metal2 38134 37145 38134 37145 0 chany_bottom_in[13]
rlabel metal1 23276 36754 23276 36754 0 chany_bottom_in[14]
rlabel metal2 9706 823 9706 823 0 chany_bottom_in[15]
rlabel via2 4922 17085 4922 17085 0 chany_bottom_in[16]
rlabel metal3 1142 7548 1142 7548 0 chany_bottom_in[17]
rlabel metal2 31602 1588 31602 1588 0 chany_bottom_in[18]
rlabel metal2 37490 1853 37490 1853 0 chany_bottom_in[1]
rlabel metal3 3902 15028 3902 15028 0 chany_bottom_in[2]
rlabel metal2 38318 7701 38318 7701 0 chany_bottom_in[3]
rlabel metal1 11362 37298 11362 37298 0 chany_bottom_in[4]
rlabel metal3 1142 38828 1142 38828 0 chany_bottom_in[5]
rlabel metal3 1142 21828 1142 21828 0 chany_bottom_in[6]
rlabel metal1 23138 1326 23138 1326 0 chany_bottom_in[7]
rlabel metal3 1142 25228 1142 25228 0 chany_bottom_in[8]
rlabel metal1 34546 37298 34546 37298 0 chany_bottom_in[9]
rlabel metal2 22586 1520 22586 1520 0 chany_bottom_out[0]
rlabel metal2 29670 1520 29670 1520 0 chany_bottom_out[10]
rlabel via2 38226 24565 38226 24565 0 chany_bottom_out[11]
rlabel metal2 38226 4913 38226 4913 0 chany_bottom_out[12]
rlabel metal1 27876 37094 27876 37094 0 chany_bottom_out[13]
rlabel metal1 37352 36346 37352 36346 0 chany_bottom_out[14]
rlabel metal1 17572 37094 17572 37094 0 chany_bottom_out[15]
rlabel metal1 1242 2822 1242 2822 0 chany_bottom_out[16]
rlabel metal2 5198 1520 5198 1520 0 chany_bottom_out[17]
rlabel metal1 14030 37094 14030 37094 0 chany_bottom_out[18]
rlabel metal1 9200 36890 9200 36890 0 chany_bottom_out[1]
rlabel metal2 38226 21233 38226 21233 0 chany_bottom_out[2]
rlabel metal2 38226 14297 38226 14297 0 chany_bottom_out[3]
rlabel metal1 38088 36890 38088 36890 0 chany_bottom_out[4]
rlabel metal2 3266 1520 3266 1520 0 chany_bottom_out[5]
rlabel metal2 38226 3077 38226 3077 0 chany_bottom_out[6]
rlabel metal2 38226 15793 38226 15793 0 chany_bottom_out[7]
rlabel metal3 1234 27268 1234 27268 0 chany_bottom_out[8]
rlabel metal1 2944 37094 2944 37094 0 chany_bottom_out[9]
rlabel metal2 36754 1588 36754 1588 0 chany_top_in[0]
rlabel metal2 2990 21199 2990 21199 0 chany_top_in[10]
rlabel metal1 828 36754 828 36754 0 chany_top_in[11]
rlabel metal1 38088 37298 38088 37298 0 chany_top_in[12]
rlabel metal2 8418 1588 8418 1588 0 chany_top_in[13]
rlabel metal2 3266 18887 3266 18887 0 chany_top_in[14]
rlabel metal2 23874 1588 23874 1588 0 chany_top_in[15]
rlabel metal2 38042 2064 38042 2064 0 chany_top_in[16]
rlabel metal1 14490 36788 14490 36788 0 chany_top_in[17]
rlabel metal2 30314 1588 30314 1588 0 chany_top_in[18]
rlabel metal2 3910 1588 3910 1588 0 chany_top_in[1]
rlabel metal3 1464 13668 1464 13668 0 chany_top_in[2]
rlabel metal2 38318 4369 38318 4369 0 chany_top_in[3]
rlabel metal2 38134 29427 38134 29427 0 chany_top_in[4]
rlabel metal1 37352 20910 37352 20910 0 chany_top_in[5]
rlabel metal2 32890 1554 32890 1554 0 chany_top_in[6]
rlabel metal3 2798 23868 2798 23868 0 chany_top_in[7]
rlabel metal1 37352 10030 37352 10030 0 chany_top_in[8]
rlabel metal3 1142 32028 1142 32028 0 chany_top_in[9]
rlabel via2 38226 22491 38226 22491 0 chany_top_out[0]
rlabel metal2 38226 34221 38226 34221 0 chany_top_out[10]
rlabel metal2 36110 1520 36110 1520 0 chany_top_out[11]
rlabel metal2 38226 36057 38226 36057 0 chany_top_out[12]
rlabel metal3 1234 33388 1234 33388 0 chany_top_out[13]
rlabel metal3 1234 2108 1234 2108 0 chany_top_out[14]
rlabel metal3 1970 12308 1970 12308 0 chany_top_out[15]
rlabel metal1 1288 2890 1288 2890 0 chany_top_out[16]
rlabel metal2 25806 1520 25806 1520 0 chany_top_out[17]
rlabel metal2 1794 37247 1794 37247 0 chany_top_out[18]
rlabel metal1 9844 37094 9844 37094 0 chany_top_out[1]
rlabel metal1 24656 37094 24656 37094 0 chany_top_out[2]
rlabel metal3 1234 29988 1234 29988 0 chany_top_out[3]
rlabel metal2 6486 1520 6486 1520 0 chany_top_out[4]
rlabel metal2 1978 1520 1978 1520 0 chany_top_out[5]
rlabel metal3 1234 8908 1234 8908 0 chany_top_out[6]
rlabel metal1 22172 36890 22172 36890 0 chany_top_out[7]
rlabel metal2 18078 1520 18078 1520 0 chany_top_out[8]
rlabel metal2 35558 37213 35558 37213 0 chany_top_out[9]
rlabel metal1 14214 17272 14214 17272 0 clknet_0_prog_clk
rlabel metal1 4600 5746 4600 5746 0 clknet_4_0_0_prog_clk
rlabel metal2 1702 17170 1702 17170 0 clknet_4_10_0_prog_clk
rlabel metal1 4002 15436 4002 15436 0 clknet_4_11_0_prog_clk
rlabel metal1 10902 12750 10902 12750 0 clknet_4_12_0_prog_clk
rlabel metal2 11730 14059 11730 14059 0 clknet_4_13_0_prog_clk
rlabel metal2 6854 17867 6854 17867 0 clknet_4_14_0_prog_clk
rlabel metal1 14950 17034 14950 17034 0 clknet_4_15_0_prog_clk
rlabel metal1 7176 5202 7176 5202 0 clknet_4_1_0_prog_clk
rlabel metal1 2346 8398 2346 8398 0 clknet_4_2_0_prog_clk
rlabel metal2 5934 6596 5934 6596 0 clknet_4_3_0_prog_clk
rlabel metal1 11868 2482 11868 2482 0 clknet_4_4_0_prog_clk
rlabel metal1 13616 5746 13616 5746 0 clknet_4_5_0_prog_clk
rlabel metal1 11914 9996 11914 9996 0 clknet_4_6_0_prog_clk
rlabel metal1 14168 11118 14168 11118 0 clknet_4_7_0_prog_clk
rlabel metal1 1656 12274 1656 12274 0 clknet_4_8_0_prog_clk
rlabel metal1 4232 12750 4232 12750 0 clknet_4_9_0_prog_clk
rlabel metal2 38318 6239 38318 6239 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal3 1740 36788 1740 36788 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 1978 8534 1978 8534 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 7222 459 7222 459 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 3818 15436 3818 15436 0 mem_bottom_track_1.DFFR_0_.D
rlabel viali 20286 3025 20286 3025 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal1 20838 5678 20838 5678 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal1 17710 1598 17710 1598 0 mem_bottom_track_1.DFFR_2_.Q
rlabel via3 7245 16524 7245 16524 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal2 13938 4760 13938 4760 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal1 13156 5814 13156 5814 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal1 9430 10098 9430 10098 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal2 23230 8636 23230 8636 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal1 10948 9010 10948 9010 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal2 21298 10353 21298 10353 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 19826 12886 19826 12886 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 8602 14382 8602 14382 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal1 1656 25874 1656 25874 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal1 1748 25806 1748 25806 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal3 7038 13260 7038 13260 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal1 1610 11050 1610 11050 0 mem_bottom_track_17.DFFR_6_.Q
rlabel metal2 2300 16560 2300 16560 0 mem_bottom_track_17.DFFR_7_.Q
rlabel metal3 2323 26316 2323 26316 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 1886 17289 1886 17289 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal2 23322 11441 23322 11441 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal1 5060 9486 5060 9486 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal1 6302 12818 6302 12818 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal2 8786 7021 8786 7021 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal1 13938 9452 13938 9452 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal1 13248 13294 13248 13294 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal2 13754 13022 13754 13022 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal1 7774 17714 7774 17714 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal1 1886 12920 1886 12920 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal1 10810 21522 10810 21522 0 mem_bottom_track_33.DFFR_5_.Q
rlabel metal3 17135 18020 17135 18020 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal1 19826 18734 19826 18734 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal1 17434 17170 17434 17170 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal1 21206 12376 21206 12376 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal1 21206 13294 21206 13294 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal1 14536 14382 14536 14382 0 mem_bottom_track_9.DFFR_5_.Q
rlabel metal2 13386 16133 13386 16133 0 mem_bottom_track_9.DFFR_6_.Q
rlabel metal1 13248 11118 13248 11118 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 16606 2414 16606 2414 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 16008 4454 16008 4454 0 mem_left_track_1.DFFR_2_.Q
rlabel metal2 13386 4182 13386 4182 0 mem_left_track_1.DFFR_3_.Q
rlabel metal1 8740 11118 8740 11118 0 mem_left_track_1.DFFR_4_.Q
rlabel metal1 9890 16592 9890 16592 0 mem_left_track_1.DFFR_5_.Q
rlabel metal2 19366 18054 19366 18054 0 mem_left_track_11.DFFR_0_.D
rlabel metal2 12558 8993 12558 8993 0 mem_left_track_11.DFFR_0_.Q
rlabel metal2 20562 4318 20562 4318 0 mem_left_track_11.DFFR_1_.Q
rlabel metal1 20608 16082 20608 16082 0 mem_left_track_13.DFFR_0_.Q
rlabel metal1 12052 14926 12052 14926 0 mem_left_track_13.DFFR_1_.Q
rlabel metal2 12052 19754 12052 19754 0 mem_left_track_15.DFFR_0_.Q
rlabel metal1 3404 18938 3404 18938 0 mem_left_track_15.DFFR_1_.Q
rlabel metal2 6256 21148 6256 21148 0 mem_left_track_17.DFFR_0_.Q
rlabel via2 6486 26333 6486 26333 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 19504 26350 19504 26350 0 mem_left_track_19.DFFR_0_.Q
rlabel via2 13846 17493 13846 17493 0 mem_left_track_19.DFFR_1_.Q
rlabel metal3 17204 13192 17204 13192 0 mem_left_track_21.DFFR_0_.Q
rlabel metal2 10902 7769 10902 7769 0 mem_left_track_21.DFFR_1_.Q
rlabel metal1 18032 18258 18032 18258 0 mem_left_track_23.DFFR_0_.Q
rlabel metal1 9016 12750 9016 12750 0 mem_left_track_23.DFFR_1_.Q
rlabel metal1 19274 15504 19274 15504 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 23874 16592 23874 16592 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 12926 16456 12926 16456 0 mem_left_track_27.DFFR_0_.Q
rlabel metal1 16560 10438 16560 10438 0 mem_left_track_27.DFFR_1_.Q
rlabel metal1 7774 4726 7774 4726 0 mem_left_track_3.DFFR_0_.Q
rlabel metal1 22494 8874 22494 8874 0 mem_left_track_3.DFFR_1_.Q
rlabel metal1 13202 2618 13202 2618 0 mem_left_track_3.DFFR_2_.Q
rlabel metal2 18354 3655 18354 3655 0 mem_left_track_3.DFFR_3_.Q
rlabel metal1 1978 12104 1978 12104 0 mem_left_track_3.DFFR_4_.Q
rlabel metal2 3450 11390 3450 11390 0 mem_left_track_3.DFFR_5_.Q
rlabel metal1 11546 21454 11546 21454 0 mem_left_track_37.DFFR_0_.Q
rlabel metal2 17250 13294 17250 13294 0 mem_left_track_5.DFFR_0_.Q
rlabel metal1 7958 21998 7958 21998 0 mem_left_track_5.DFFR_1_.Q
rlabel metal1 5106 4046 5106 4046 0 mem_left_track_5.DFFR_2_.Q
rlabel metal1 6348 7786 6348 7786 0 mem_left_track_5.DFFR_3_.Q
rlabel metal1 7314 10098 7314 10098 0 mem_left_track_5.DFFR_4_.Q
rlabel metal1 19458 12784 19458 12784 0 mem_left_track_5.DFFR_5_.Q
rlabel metal1 5927 16762 5927 16762 0 mem_left_track_7.DFFR_0_.Q
rlabel metal1 7636 16422 7636 16422 0 mem_left_track_7.DFFR_1_.Q
rlabel metal2 5750 18734 5750 18734 0 mem_left_track_7.DFFR_2_.Q
rlabel metal1 5980 18190 5980 18190 0 mem_left_track_7.DFFR_3_.Q
rlabel metal1 1886 16626 1886 16626 0 mem_left_track_7.DFFR_4_.Q
rlabel metal1 3174 16422 3174 16422 0 mem_left_track_7.DFFR_5_.Q
rlabel metal2 21942 16286 21942 16286 0 mem_left_track_9.DFFR_0_.Q
rlabel metal2 7130 18615 7130 18615 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 8326 17102 8326 17102 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 20562 13396 20562 13396 0 mem_top_track_0.DFFR_2_.Q
rlabel metal1 12788 21046 12788 21046 0 mem_top_track_0.DFFR_3_.Q
rlabel metal1 8671 19278 8671 19278 0 mem_top_track_0.DFFR_4_.Q
rlabel metal1 10327 14994 10327 14994 0 mem_top_track_0.DFFR_5_.Q
rlabel metal1 1886 15096 1886 15096 0 mem_top_track_0.DFFR_6_.Q
rlabel metal2 16146 15181 16146 15181 0 mem_top_track_0.DFFR_7_.Q
rlabel metal1 8924 3910 8924 3910 0 mem_top_track_16.DFFR_0_.D
rlabel metal2 22034 14722 22034 14722 0 mem_top_track_16.DFFR_0_.Q
rlabel metal2 2392 17476 2392 17476 0 mem_top_track_16.DFFR_1_.Q
rlabel metal1 4876 14382 4876 14382 0 mem_top_track_16.DFFR_2_.Q
rlabel metal1 16054 19822 16054 19822 0 mem_top_track_16.DFFR_3_.Q
rlabel metal1 1971 6970 1971 6970 0 mem_top_track_16.DFFR_4_.Q
rlabel metal1 1978 5576 1978 5576 0 mem_top_track_16.DFFR_5_.Q
rlabel via2 19642 3043 19642 3043 0 mem_top_track_16.DFFR_6_.Q
rlabel metal2 14306 6681 14306 6681 0 mem_top_track_16.DFFR_7_.Q
rlabel metal2 12466 23936 12466 23936 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 9062 25262 9062 25262 0 mem_top_track_24.DFFR_1_.Q
rlabel metal2 5750 16473 5750 16473 0 mem_top_track_24.DFFR_2_.Q
rlabel metal1 13984 27438 13984 27438 0 mem_top_track_24.DFFR_3_.Q
rlabel metal1 5934 15606 5934 15606 0 mem_top_track_24.DFFR_4_.Q
rlabel metal1 11500 20910 11500 20910 0 mem_top_track_24.DFFR_5_.Q
rlabel metal1 9246 13226 9246 13226 0 mem_top_track_24.DFFR_6_.Q
rlabel metal1 14582 14552 14582 14552 0 mem_top_track_24.DFFR_7_.Q
rlabel metal2 14490 27166 14490 27166 0 mem_top_track_32.DFFR_0_.Q
rlabel metal2 9430 14076 9430 14076 0 mem_top_track_32.DFFR_1_.Q
rlabel metal2 1978 17340 1978 17340 0 mem_top_track_32.DFFR_2_.Q
rlabel metal1 3266 17782 3266 17782 0 mem_top_track_32.DFFR_3_.Q
rlabel metal2 13662 17255 13662 17255 0 mem_top_track_32.DFFR_4_.Q
rlabel metal1 16560 15402 16560 15402 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 20056 13226 20056 13226 0 mem_top_track_8.DFFR_1_.Q
rlabel metal1 17158 17714 17158 17714 0 mem_top_track_8.DFFR_2_.Q
rlabel metal1 15042 6086 15042 6086 0 mem_top_track_8.DFFR_3_.Q
rlabel metal1 6486 4046 6486 4046 0 mem_top_track_8.DFFR_4_.Q
rlabel metal1 14766 7752 14766 7752 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 21298 8874 21298 8874 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 20700 9486 20700 9486 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal2 21758 4675 21758 4675 0 mux_bottom_track_1.INVTX1_3_.out
rlabel via1 20102 3621 20102 3621 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal1 17710 13838 17710 13838 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal1 18676 18326 18676 18326 0 mux_bottom_track_1.INVTX1_6_.out
rlabel metal1 8832 21454 8832 21454 0 mux_bottom_track_1.INVTX1_7_.out
rlabel metal1 17342 20978 17342 20978 0 mux_bottom_track_1.INVTX1_8_.out
rlabel metal1 20884 7242 20884 7242 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 18262 5712 18262 5712 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 18308 9962 18308 9962 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 21597 3026 21597 3026 0 mux_bottom_track_1.out
rlabel metal2 16974 8942 16974 8942 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 7544 25806 7544 25806 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal2 19734 13770 19734 13770 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 2254 21454 2254 21454 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal2 21114 10132 21114 10132 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 20884 11662 20884 11662 0 mux_bottom_track_17.INVTX1_5_.out
rlabel metal2 10672 22080 10672 22080 0 mux_bottom_track_17.INVTX1_6_.out
rlabel metal1 29371 11526 29371 11526 0 mux_bottom_track_17.INVTX1_7_.out
rlabel metal3 16537 20740 16537 20740 0 mux_bottom_track_17.INVTX1_8_.out
rlabel metal3 17687 20876 17687 20876 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel via2 12742 19669 12742 19669 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 4922 21386 4922 21386 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 2760 19686 2760 19686 0 mux_bottom_track_17.out
rlabel metal1 13110 23188 13110 23188 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal2 13754 24514 13754 24514 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal1 15410 20332 15410 20332 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal2 1794 19789 1794 19789 0 mux_bottom_track_25.INVTX1_3_.out
rlabel metal1 2944 22678 2944 22678 0 mux_bottom_track_25.INVTX1_4_.out
rlabel metal1 14398 20808 14398 20808 0 mux_bottom_track_25.INVTX1_5_.out
rlabel metal1 21804 4454 21804 4454 0 mux_bottom_track_25.INVTX1_6_.out
rlabel metal2 19458 4811 19458 4811 0 mux_bottom_track_25.INVTX1_7_.out
rlabel via2 15686 20349 15686 20349 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 14674 17408 14674 17408 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 18170 8398 18170 8398 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 32361 8466 32361 8466 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 35098 7854 35098 7854 0 mux_bottom_track_25.out
rlabel metal1 23138 21386 23138 21386 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal1 19734 23630 19734 23630 0 mux_bottom_track_33.INVTX1_1_.out
rlabel metal2 32430 24072 32430 24072 0 mux_bottom_track_33.INVTX1_2_.out
rlabel metal1 9614 24106 9614 24106 0 mux_bottom_track_33.INVTX1_3_.out
rlabel metal2 9246 22219 9246 22219 0 mux_bottom_track_33.INVTX1_4_.out
rlabel metal1 25116 16626 25116 16626 0 mux_bottom_track_33.INVTX1_5_.out
rlabel metal2 17158 27948 17158 27948 0 mux_bottom_track_33.INVTX1_6_.out
rlabel metal1 10718 21046 10718 21046 0 mux_bottom_track_33.INVTX1_7_.out
rlabel metal2 20378 20570 20378 20570 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 21666 19856 21666 19856 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 17618 24888 17618 24888 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 13156 19754 13156 19754 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 3450 6290 3450 6290 0 mux_bottom_track_33.out
rlabel metal1 17434 8874 17434 8874 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 20332 14926 20332 14926 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal2 18630 14892 18630 14892 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal1 14720 2822 14720 2822 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal1 21068 31926 21068 31926 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal1 16560 24582 16560 24582 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal1 14306 18666 14306 18666 0 mux_bottom_track_9.INVTX1_6_.out
rlabel metal2 12558 24735 12558 24735 0 mux_bottom_track_9.INVTX1_7_.out
rlabel metal1 18906 20366 18906 20366 0 mux_bottom_track_9.INVTX1_8_.out
rlabel metal1 19228 14314 19228 14314 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 15916 18802 15916 18802 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 35558 28016 35558 28016 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36202 36550 36202 36550 0 mux_bottom_track_9.out
rlabel via2 19366 6749 19366 6749 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 20930 12614 20930 12614 0 mux_left_track_1.INVTX1_2_.out
rlabel via2 2162 23613 2162 23613 0 mux_left_track_1.INVTX1_3_.out
rlabel metal1 17342 8942 17342 8942 0 mux_left_track_1.INVTX1_4_.out
rlabel metal2 16606 11764 16606 11764 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal2 15226 7072 15226 7072 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 17434 11050 17434 11050 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 2254 24752 2254 24752 0 mux_left_track_1.out
rlabel metal1 16928 19686 16928 19686 0 mux_left_track_11.INVTX1_1_.out
rlabel metal2 28198 5287 28198 5287 0 mux_left_track_11.INVTX1_2_.out
rlabel metal1 15778 5134 15778 5134 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21942 6630 21942 6630 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 16560 5202 16560 5202 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 28014 3553 28014 3553 0 mux_left_track_11.out
rlabel metal1 17710 16014 17710 16014 0 mux_left_track_13.INVTX1_1_.out
rlabel metal1 20424 15062 20424 15062 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 26818 16048 26818 16048 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 33120 17170 33120 17170 0 mux_left_track_13.out
rlabel metal1 15226 26452 15226 26452 0 mux_left_track_15.INVTX1_1_.out
rlabel metal2 8326 24922 8326 24922 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 4462 23562 4462 23562 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 5934 28118 5934 28118 0 mux_left_track_15.out
rlabel metal1 13708 26894 13708 26894 0 mux_left_track_17.INVTX1_1_.out
rlabel metal1 11132 26486 11132 26486 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9154 27030 9154 27030 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5750 31790 5750 31790 0 mux_left_track_17.out
rlabel metal1 18354 27846 18354 27846 0 mux_left_track_19.INVTX1_1_.out
rlabel metal1 19228 23834 19228 23834 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 21988 25126 21988 25126 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 20930 24480 20930 24480 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 31786 28356 31786 28356 0 mux_left_track_19.out
rlabel metal1 22632 16422 22632 16422 0 mux_left_track_21.INVTX1_1_.out
rlabel metal1 23046 8364 23046 8364 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 24518 9996 24518 9996 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25714 8398 25714 8398 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 26174 7310 26174 7310 0 mux_left_track_21.out
rlabel metal1 20608 17714 20608 17714 0 mux_left_track_23.INVTX1_1_.out
rlabel metal1 16882 10676 16882 10676 0 mux_left_track_23.INVTX1_2_.out
rlabel metal2 21482 16014 21482 16014 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 26818 14144 26818 14144 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 26634 14144 26634 14144 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30912 13906 30912 13906 0 mux_left_track_23.out
rlabel metal2 21850 15266 21850 15266 0 mux_left_track_25.INVTX1_1_.out
rlabel metal2 16974 20706 16974 20706 0 mux_left_track_25.INVTX1_2_.out
rlabel metal1 22770 15674 22770 15674 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22402 20944 22402 20944 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23874 21046 23874 21046 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 29900 25262 29900 25262 0 mux_left_track_25.out
rlabel metal1 12650 22542 12650 22542 0 mux_left_track_27.INVTX1_1_.out
rlabel metal1 13524 19278 13524 19278 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 29854 4794 29854 4794 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel viali 30958 4588 30958 4588 0 mux_left_track_27.out
rlabel metal1 20562 7922 20562 7922 0 mux_left_track_3.INVTX1_1_.out
rlabel metal2 17158 7531 17158 7531 0 mux_left_track_3.INVTX1_2_.out
rlabel metal2 17526 8704 17526 8704 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal2 19826 8160 19826 8160 0 mux_left_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 6164 19754 6164 19754 0 mux_left_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 7590 31450 7590 31450 0 mux_left_track_3.out
rlabel metal1 3312 20366 3312 20366 0 mux_left_track_37.INVTX1_0_.out
rlabel metal2 11454 21267 11454 21267 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 26680 20366 26680 20366 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 34914 18258 34914 18258 0 mux_left_track_37.out
rlabel metal1 7406 20842 7406 20842 0 mux_left_track_5.INVTX1_1_.out
rlabel metal1 15916 3570 15916 3570 0 mux_left_track_5.INVTX1_2_.out
rlabel metal1 16560 12138 16560 12138 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel via3 14283 13668 14283 13668 0 mux_left_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 21712 16660 21712 16660 0 mux_left_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 32798 20876 32798 20876 0 mux_left_track_5.out
rlabel metal2 5934 20604 5934 20604 0 mux_left_track_7.INVTX1_1_.out
rlabel metal1 15088 31858 15088 31858 0 mux_left_track_7.INVTX1_2_.out
rlabel metal1 8004 24718 8004 24718 0 mux_left_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 7544 21964 7544 21964 0 mux_left_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 14168 34578 14168 34578 0 mux_left_track_7.out
rlabel metal1 8418 22712 8418 22712 0 mux_left_track_9.INVTX1_1_.out
rlabel via3 20171 8772 20171 8772 0 mux_left_track_9.INVTX1_2_.out
rlabel via1 23414 21522 23414 21522 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 22954 18666 22954 18666 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23874 18802 23874 18802 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30958 28050 30958 28050 0 mux_left_track_9.out
rlabel metal1 27186 22066 27186 22066 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 9154 31926 9154 31926 0 mux_top_track_0.INVTX1_1_.out
rlabel metal2 19550 20060 19550 20060 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 25714 16218 25714 16218 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 15088 15062 15088 15062 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 38042 22202 38042 22202 0 mux_top_track_0.out
rlabel metal1 21068 31994 21068 31994 0 mux_top_track_16.INVTX1_0_.out
rlabel metal1 1840 26758 1840 26758 0 mux_top_track_16.INVTX1_1_.out
rlabel metal1 2668 20502 2668 20502 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 14766 12614 14766 12614 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 18676 4046 18676 4046 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 23506 2992 23506 2992 0 mux_top_track_16.out
rlabel metal1 20838 32742 20838 32742 0 mux_top_track_24.INVTX1_0_.out
rlabel metal2 8602 27166 8602 27166 0 mux_top_track_24.INVTX1_1_.out
rlabel metal1 13202 23596 13202 23596 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 13754 21386 13754 21386 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 36018 30566 36018 30566 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 36432 34714 36432 34714 0 mux_top_track_24.out
rlabel metal1 6256 32742 6256 32742 0 mux_top_track_32.INVTX1_0_.out
rlabel metal2 21482 19618 21482 19618 0 mux_top_track_32.INVTX1_1_.out
rlabel metal2 6946 20162 6946 20162 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 17986 25772 17986 25772 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15134 21046 15134 21046 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 15410 17527 15410 17527 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel via2 1978 6307 1978 6307 0 mux_top_track_32.out
rlabel metal2 22770 2737 22770 2737 0 mux_top_track_8.INVTX1_0_.out
rlabel metal1 24794 3094 24794 3094 0 mux_top_track_8.INVTX1_1_.out
rlabel metal2 17802 5015 17802 5015 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20378 17544 20378 17544 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19688 4794 19688 4794 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 19090 6256 19090 6256 0 mux_top_track_8.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 27370 3468 27370 3468 0 mux_top_track_8.out
rlabel metal2 2714 25503 2714 25503 0 net1
rlabel metal2 33074 9622 33074 9622 0 net10
rlabel metal1 3128 31790 3128 31790 0 net100
rlabel metal1 4600 31994 4600 31994 0 net101
rlabel metal2 33258 30838 33258 30838 0 net102
rlabel metal1 22678 2448 22678 2448 0 net103
rlabel metal2 13110 23936 13110 23936 0 net104
rlabel metal2 34546 24038 34546 24038 0 net105
rlabel metal2 38042 6460 38042 6460 0 net106
rlabel metal2 27830 37060 27830 37060 0 net107
rlabel metal2 37306 35666 37306 35666 0 net108
rlabel metal2 17526 34485 17526 34485 0 net109
rlabel metal1 3818 7208 3818 7208 0 net11
rlabel metal2 2438 4590 2438 4590 0 net110
rlabel metal2 5290 2125 5290 2125 0 net111
rlabel metal1 13754 36890 13754 36890 0 net112
rlabel metal2 9154 36550 9154 36550 0 net113
rlabel metal2 38042 20196 38042 20196 0 net114
rlabel metal2 37306 13804 37306 13804 0 net115
rlabel metal1 36662 36720 36662 36720 0 net116
rlabel via3 3197 2652 3197 2652 0 net117
rlabel metal1 37996 3502 37996 3502 0 net118
rlabel metal2 36570 15334 36570 15334 0 net119
rlabel metal3 4508 19380 4508 19380 0 net12
rlabel metal1 1610 27404 1610 27404 0 net120
rlabel metal2 20746 21794 20746 21794 0 net121
rlabel metal2 37858 22406 37858 22406 0 net122
rlabel metal1 38042 34612 38042 34612 0 net123
rlabel metal1 36041 2414 36041 2414 0 net124
rlabel metal1 38042 36176 38042 36176 0 net125
rlabel metal1 4255 33490 4255 33490 0 net126
rlabel metal2 21298 15385 21298 15385 0 net127
rlabel metal2 13754 18173 13754 18173 0 net128
rlabel metal2 2346 4556 2346 4556 0 net129
rlabel metal1 24656 30702 24656 30702 0 net13
rlabel metal1 25944 9894 25944 9894 0 net130
rlabel metal3 2047 35972 2047 35972 0 net131
rlabel metal1 9660 37298 9660 37298 0 net132
rlabel metal1 23000 34510 23000 34510 0 net133
rlabel metal1 6348 23834 6348 23834 0 net134
rlabel metal2 6578 2193 6578 2193 0 net135
rlabel metal1 3772 2550 3772 2550 0 net136
rlabel metal2 1564 16626 1564 16626 0 net137
rlabel metal1 20056 36754 20056 36754 0 net138
rlabel metal1 18170 2380 18170 2380 0 net139
rlabel metal2 4094 24786 4094 24786 0 net14
rlabel metal1 36110 37230 36110 37230 0 net140
rlabel metal2 14858 1010 14858 1010 0 net141
rlabel metal1 16560 14926 16560 14926 0 net142
rlabel metal2 13570 8296 13570 8296 0 net143
rlabel metal2 13570 20196 13570 20196 0 net144
rlabel metal2 22678 8466 22678 8466 0 net145
rlabel metal1 18998 16014 18998 16014 0 net146
rlabel metal1 2507 20978 2507 20978 0 net147
rlabel metal1 19274 4012 19274 4012 0 net148
rlabel metal1 13754 22712 13754 22712 0 net149
rlabel metal1 12696 37094 12696 37094 0 net15
rlabel metal1 19734 10098 19734 10098 0 net150
rlabel metal2 16974 24922 16974 24922 0 net151
rlabel metal1 10166 19890 10166 19890 0 net152
rlabel metal1 4186 14484 4186 14484 0 net153
rlabel metal1 18630 11662 18630 11662 0 net154
rlabel metal2 6762 24990 6762 24990 0 net155
rlabel metal2 24978 19040 24978 19040 0 net156
rlabel metal2 23414 7072 23414 7072 0 net157
rlabel metal1 21068 25262 21068 25262 0 net158
rlabel metal1 26220 10574 26220 10574 0 net159
rlabel metal2 38134 11526 38134 11526 0 net16
rlabel metal2 26726 14688 26726 14688 0 net160
rlabel metal1 21896 21522 21896 21522 0 net161
rlabel metal2 24610 15776 24610 15776 0 net162
rlabel metal1 3496 21454 3496 21454 0 net163
rlabel metal1 8648 24242 8648 24242 0 net164
rlabel metal1 23736 10098 23736 10098 0 net165
rlabel metal1 25300 20366 25300 20366 0 net166
rlabel metal1 27232 6222 27232 6222 0 net17
rlabel metal1 4646 37128 4646 37128 0 net18
rlabel metal1 34270 36550 34270 36550 0 net19
rlabel metal2 5842 34748 5842 34748 0 net2
rlabel metal2 37490 33116 37490 33116 0 net20
rlabel metal1 24840 5678 24840 5678 0 net21
rlabel metal1 20102 2550 20102 2550 0 net22
rlabel metal2 36018 25469 36018 25469 0 net23
rlabel metal2 38134 12410 38134 12410 0 net24
rlabel metal1 15364 28526 15364 28526 0 net25
rlabel metal2 30774 6052 30774 6052 0 net26
rlabel metal2 33074 33694 33074 33694 0 net27
rlabel metal2 23414 2329 23414 2329 0 net28
rlabel metal1 6578 29682 6578 29682 0 net29
rlabel metal1 13156 1190 13156 1190 0 net3
rlabel metal1 21965 4590 21965 4590 0 net30
rlabel metal1 37053 3910 37053 3910 0 net31
rlabel metal1 20562 37162 20562 37162 0 net32
rlabel metal1 19412 37094 19412 37094 0 net33
rlabel metal1 20792 36822 20792 36822 0 net34
rlabel metal1 38088 36550 38088 36550 0 net35
rlabel metal1 22126 36686 22126 36686 0 net36
rlabel metal1 20286 3502 20286 3502 0 net37
rlabel metal2 6762 17017 6762 17017 0 net38
rlabel metal1 2530 10676 2530 10676 0 net39
rlabel metal1 20654 2856 20654 2856 0 net4
rlabel metal2 32338 3672 32338 3672 0 net40
rlabel metal2 37766 3366 37766 3366 0 net41
rlabel metal1 6900 14858 6900 14858 0 net42
rlabel metal1 34937 7990 34937 7990 0 net43
rlabel metal1 11914 37230 11914 37230 0 net44
rlabel metal1 5244 37230 5244 37230 0 net45
rlabel metal2 4002 21828 4002 21828 0 net46
rlabel metal1 16744 5678 16744 5678 0 net47
rlabel metal1 17986 25840 17986 25840 0 net48
rlabel metal1 35328 37230 35328 37230 0 net49
rlabel metal2 5198 25806 5198 25806 0 net5
rlabel metal2 37766 2108 37766 2108 0 net50
rlabel metal2 14858 23460 14858 23460 0 net51
rlabel metal2 1886 33660 1886 33660 0 net52
rlabel metal1 37766 37196 37766 37196 0 net53
rlabel metal1 9338 2482 9338 2482 0 net54
rlabel metal2 18492 18836 18492 18836 0 net55
rlabel metal1 24472 2618 24472 2618 0 net56
rlabel metal1 36731 3638 36731 3638 0 net57
rlabel metal1 13846 36754 13846 36754 0 net58
rlabel metal1 31510 21522 31510 21522 0 net59
rlabel metal2 2898 7905 2898 7905 0 net6
rlabel metal1 10258 2346 10258 2346 0 net60
rlabel metal1 16928 12750 16928 12750 0 net61
rlabel metal2 34086 5542 34086 5542 0 net62
rlabel metal1 37996 29478 37996 29478 0 net63
rlabel metal1 37812 20910 37812 20910 0 net64
rlabel metal1 33810 9962 33810 9962 0 net65
rlabel metal1 4462 24174 4462 24174 0 net66
rlabel metal2 34546 12342 34546 12342 0 net67
rlabel metal1 5612 32334 5612 32334 0 net68
rlabel metal2 38134 8500 38134 8500 0 net69
rlabel metal2 37030 28764 37030 28764 0 net7
rlabel metal1 4600 36006 4600 36006 0 net70
rlabel metal1 1656 23698 1656 23698 0 net71
rlabel metal2 20102 2176 20102 2176 0 net72
rlabel metal2 16514 8058 16514 8058 0 net73
rlabel metal2 34638 25092 34638 25092 0 net74
rlabel metal1 22356 2618 22356 2618 0 net75
rlabel metal1 29210 37094 29210 37094 0 net76
rlabel metal1 26174 32878 26174 32878 0 net77
rlabel metal1 4324 36550 4324 36550 0 net78
rlabel metal2 6578 34476 6578 34476 0 net79
rlabel metal2 21390 3332 21390 3332 0 net8
rlabel metal1 26266 2618 26266 2618 0 net80
rlabel metal3 2277 26588 2277 26588 0 net81
rlabel metal1 2852 34918 2852 34918 0 net82
rlabel metal1 37007 19482 37007 19482 0 net83
rlabel metal2 37766 21777 37766 21777 0 net84
rlabel metal1 2392 23494 2392 23494 0 net85
rlabel metal1 25438 2414 25438 2414 0 net86
rlabel metal2 34822 13668 34822 13668 0 net87
rlabel metal1 36984 27438 36984 27438 0 net88
rlabel metal1 34684 2414 34684 2414 0 net89
rlabel metal1 23552 31858 23552 31858 0 net9
rlabel metal2 32338 29444 32338 29444 0 net90
rlabel metal2 20102 30804 20102 30804 0 net91
rlabel metal2 33718 16524 33718 16524 0 net92
rlabel metal2 38042 17306 38042 17306 0 net93
rlabel metal1 7682 31994 7682 31994 0 net94
rlabel metal2 36110 22644 36110 22644 0 net95
rlabel metal1 16146 36754 16146 36754 0 net96
rlabel metal2 36478 30532 36478 30532 0 net97
rlabel metal2 1610 3723 1610 3723 0 net98
rlabel metal1 34868 17306 34868 17306 0 net99
rlabel metal2 14214 2251 14214 2251 0 pReset
rlabel metal2 4094 3587 4094 3587 0 prog_clk
rlabel metal3 38786 25908 38786 25908 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 21942 1588 21942 1588 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal1 29808 37230 29808 37230 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 28566 37230 28566 37230 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 3082 36788 3082 36788 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 6624 37230 6624 37230 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 27094 1588 27094 1588 0 top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 2806 9605 2806 9605 0 top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal3 1234 34748 1234 34748 0 top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 38318 19227 38318 19227 0 top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
