magic
tech sky130A
magscale 1 2
timestamp 1672417964
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 14 1368 29978 27792
<< metal2 >>
rect 662 29200 718 29800
rect 1950 29200 2006 29800
rect 3238 29200 3294 29800
rect 3882 29200 3938 29800
rect 5170 29200 5226 29800
rect 6458 29200 6514 29800
rect 7746 29200 7802 29800
rect 9034 29200 9090 29800
rect 10322 29200 10378 29800
rect 10966 29200 11022 29800
rect 12254 29200 12310 29800
rect 13542 29200 13598 29800
rect 14830 29200 14886 29800
rect 16118 29200 16174 29800
rect 16762 29200 16818 29800
rect 18050 29200 18106 29800
rect 19338 29200 19394 29800
rect 20626 29200 20682 29800
rect 21914 29200 21970 29800
rect 23202 29200 23258 29800
rect 23846 29200 23902 29800
rect 25134 29200 25190 29800
rect 26422 29200 26478 29800
rect 27710 29200 27766 29800
rect 28998 29200 29054 29800
rect 29642 29200 29698 29800
rect 18 200 74 800
rect 662 200 718 800
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 6458 200 6514 800
rect 7746 200 7802 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 17406 200 17462 800
rect 18694 200 18750 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 21914 200 21970 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 28998 200 29054 800
<< obsm2 >>
rect 20 29144 606 29345
rect 774 29144 1894 29345
rect 2062 29144 3182 29345
rect 3350 29144 3826 29345
rect 3994 29144 5114 29345
rect 5282 29144 6402 29345
rect 6570 29144 7690 29345
rect 7858 29144 8978 29345
rect 9146 29144 10266 29345
rect 10434 29144 10910 29345
rect 11078 29144 12198 29345
rect 12366 29144 13486 29345
rect 13654 29144 14774 29345
rect 14942 29144 16062 29345
rect 16230 29144 16706 29345
rect 16874 29144 17994 29345
rect 18162 29144 19282 29345
rect 19450 29144 20570 29345
rect 20738 29144 21858 29345
rect 22026 29144 23146 29345
rect 23314 29144 23790 29345
rect 23958 29144 25078 29345
rect 25246 29144 26366 29345
rect 26534 29144 27654 29345
rect 27822 29144 28942 29345
rect 29110 29144 29586 29345
rect 29754 29144 29974 29345
rect 20 856 29974 29144
rect 130 144 606 856
rect 774 144 1894 856
rect 2062 144 3182 856
rect 3350 144 4470 856
rect 4638 144 5758 856
rect 5926 144 6402 856
rect 6570 144 7690 856
rect 7858 144 8978 856
rect 9146 144 10266 856
rect 10434 144 11554 856
rect 11722 144 12842 856
rect 13010 144 13486 856
rect 13654 144 14774 856
rect 14942 144 16062 856
rect 16230 144 17350 856
rect 17518 144 18638 856
rect 18806 144 19282 856
rect 19450 144 20570 856
rect 20738 144 21858 856
rect 22026 144 23146 856
rect 23314 144 24434 856
rect 24602 144 25722 856
rect 25890 144 26366 856
rect 26534 144 27654 856
rect 27822 144 28942 856
rect 29110 144 29974 856
rect 20 31 29974 144
<< metal3 >>
rect 200 29248 800 29368
rect 29200 28568 29800 28688
rect 200 27888 800 28008
rect 200 27208 800 27328
rect 29200 27208 29800 27328
rect 200 25848 800 25968
rect 29200 25848 29800 25968
rect 200 24488 800 24608
rect 29200 24488 29800 24608
rect 200 23128 800 23248
rect 29200 23128 29800 23248
rect 29200 22448 29800 22568
rect 200 21768 800 21888
rect 29200 21088 29800 21208
rect 200 20408 800 20528
rect 200 19728 800 19848
rect 29200 19728 29800 19848
rect 200 18368 800 18488
rect 29200 18368 29800 18488
rect 200 17008 800 17128
rect 29200 17008 29800 17128
rect 200 15648 800 15768
rect 29200 15648 29800 15768
rect 29200 14968 29800 15088
rect 200 14288 800 14408
rect 200 13608 800 13728
rect 29200 13608 29800 13728
rect 200 12248 800 12368
rect 29200 12248 29800 12368
rect 200 10888 800 11008
rect 29200 10888 29800 11008
rect 200 9528 800 9648
rect 29200 9528 29800 9648
rect 29200 8848 29800 8968
rect 200 8168 800 8288
rect 29200 7488 29800 7608
rect 200 6808 800 6928
rect 200 6128 800 6248
rect 29200 6128 29800 6248
rect 200 4768 800 4888
rect 29200 4768 29800 4888
rect 200 3408 800 3528
rect 29200 3408 29800 3528
rect 200 2048 800 2168
rect 29200 2048 29800 2168
rect 29200 1368 29800 1488
rect 200 688 800 808
rect 29200 8 29800 128
<< obsm3 >>
rect 880 29168 29979 29341
rect 800 28768 29979 29168
rect 800 28488 29120 28768
rect 29880 28488 29979 28768
rect 800 28088 29979 28488
rect 880 27808 29979 28088
rect 800 27408 29979 27808
rect 880 27128 29120 27408
rect 29880 27128 29979 27408
rect 800 26048 29979 27128
rect 880 25768 29120 26048
rect 29880 25768 29979 26048
rect 800 24688 29979 25768
rect 880 24408 29120 24688
rect 29880 24408 29979 24688
rect 800 23328 29979 24408
rect 880 23048 29120 23328
rect 29880 23048 29979 23328
rect 800 22648 29979 23048
rect 800 22368 29120 22648
rect 29880 22368 29979 22648
rect 800 21968 29979 22368
rect 880 21688 29979 21968
rect 800 21288 29979 21688
rect 800 21008 29120 21288
rect 29880 21008 29979 21288
rect 800 20608 29979 21008
rect 880 20328 29979 20608
rect 800 19928 29979 20328
rect 880 19648 29120 19928
rect 29880 19648 29979 19928
rect 800 18568 29979 19648
rect 880 18288 29120 18568
rect 29880 18288 29979 18568
rect 800 17208 29979 18288
rect 880 16928 29120 17208
rect 29880 16928 29979 17208
rect 800 15848 29979 16928
rect 880 15568 29120 15848
rect 29880 15568 29979 15848
rect 800 15168 29979 15568
rect 800 14888 29120 15168
rect 29880 14888 29979 15168
rect 800 14488 29979 14888
rect 880 14208 29979 14488
rect 800 13808 29979 14208
rect 880 13528 29120 13808
rect 29880 13528 29979 13808
rect 800 12448 29979 13528
rect 880 12168 29120 12448
rect 29880 12168 29979 12448
rect 800 11088 29979 12168
rect 880 10808 29120 11088
rect 29880 10808 29979 11088
rect 800 9728 29979 10808
rect 880 9448 29120 9728
rect 29880 9448 29979 9728
rect 800 9048 29979 9448
rect 800 8768 29120 9048
rect 29880 8768 29979 9048
rect 800 8368 29979 8768
rect 880 8088 29979 8368
rect 800 7688 29979 8088
rect 800 7408 29120 7688
rect 29880 7408 29979 7688
rect 800 7008 29979 7408
rect 880 6728 29979 7008
rect 800 6328 29979 6728
rect 880 6048 29120 6328
rect 29880 6048 29979 6328
rect 800 4968 29979 6048
rect 880 4688 29120 4968
rect 29880 4688 29979 4968
rect 800 3608 29979 4688
rect 880 3328 29120 3608
rect 29880 3328 29979 3608
rect 800 2248 29979 3328
rect 880 1968 29120 2248
rect 29880 1968 29979 2248
rect 800 1568 29979 1968
rect 800 1288 29120 1568
rect 29880 1288 29979 1568
rect 800 888 29979 1288
rect 880 608 29979 888
rect 800 208 29979 608
rect 800 35 29120 208
rect 29880 35 29979 208
<< metal4 >>
rect 4417 2128 4737 27792
rect 7890 2128 8210 27792
rect 11363 2128 11683 27792
rect 14836 2128 15156 27792
rect 18309 2128 18629 27792
rect 21782 2128 22102 27792
rect 25255 2128 25575 27792
rect 28728 2128 29048 27792
<< obsm4 >>
rect 12939 3027 14756 25397
rect 15236 3027 18229 25397
rect 18709 3027 21702 25397
rect 22182 3027 23861 25397
<< labels >>
rlabel metal2 s 5170 29200 5226 29800 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 1 nsew signal input
rlabel metal2 s 3238 29200 3294 29800 6 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 2 nsew signal input
rlabel metal3 s 200 20408 800 20528 6 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 3 nsew signal input
rlabel metal3 s 29200 8848 29800 8968 6 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 4 nsew signal input
rlabel metal3 s 29200 18368 29800 18488 6 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 5 nsew signal input
rlabel metal2 s 16762 29200 16818 29800 6 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 6 nsew signal input
rlabel metal2 s 7746 200 7802 800 6 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 7 nsew signal input
rlabel metal2 s 11610 200 11666 800 6 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 8 nsew signal input
rlabel metal2 s 24490 200 24546 800 6 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 9 nsew signal input
rlabel metal3 s 200 688 800 808 6 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 10 nsew signal input
rlabel metal3 s 29200 23128 29800 23248 6 ccff_head
port 11 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 ccff_tail
port 12 nsew signal output
rlabel metal2 s 25778 200 25834 800 6 chanx_left_in[0]
port 13 nsew signal input
rlabel metal3 s 200 24488 800 24608 6 chanx_left_in[10]
port 14 nsew signal input
rlabel metal2 s 25134 29200 25190 29800 6 chanx_left_in[11]
port 15 nsew signal input
rlabel metal3 s 29200 14968 29800 15088 6 chanx_left_in[12]
port 16 nsew signal input
rlabel metal2 s 9034 29200 9090 29800 6 chanx_left_in[13]
port 17 nsew signal input
rlabel metal3 s 200 27888 800 28008 6 chanx_left_in[14]
port 18 nsew signal input
rlabel metal3 s 200 19728 800 19848 6 chanx_left_in[15]
port 19 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 chanx_left_in[16]
port 20 nsew signal input
rlabel metal3 s 200 13608 800 13728 6 chanx_left_in[17]
port 21 nsew signal input
rlabel metal3 s 29200 25848 29800 25968 6 chanx_left_in[18]
port 22 nsew signal input
rlabel metal3 s 29200 3408 29800 3528 6 chanx_left_in[1]
port 23 nsew signal input
rlabel metal2 s 19338 29200 19394 29800 6 chanx_left_in[2]
port 24 nsew signal input
rlabel metal3 s 200 15648 800 15768 6 chanx_left_in[3]
port 25 nsew signal input
rlabel metal2 s 10966 29200 11022 29800 6 chanx_left_in[4]
port 26 nsew signal input
rlabel metal2 s 12254 29200 12310 29800 6 chanx_left_in[5]
port 27 nsew signal input
rlabel metal2 s 21914 29200 21970 29800 6 chanx_left_in[6]
port 28 nsew signal input
rlabel metal3 s 200 21768 800 21888 6 chanx_left_in[7]
port 29 nsew signal input
rlabel metal3 s 29200 28568 29800 28688 6 chanx_left_in[8]
port 30 nsew signal input
rlabel metal3 s 29200 24488 29800 24608 6 chanx_left_in[9]
port 31 nsew signal input
rlabel metal3 s 29200 27208 29800 27328 6 chanx_left_out[0]
port 32 nsew signal output
rlabel metal3 s 29200 6128 29800 6248 6 chanx_left_out[10]
port 33 nsew signal output
rlabel metal2 s 18050 29200 18106 29800 6 chanx_left_out[11]
port 34 nsew signal output
rlabel metal2 s 13542 29200 13598 29800 6 chanx_left_out[12]
port 35 nsew signal output
rlabel metal3 s 200 3408 800 3528 6 chanx_left_out[13]
port 36 nsew signal output
rlabel metal3 s 200 29248 800 29368 6 chanx_left_out[14]
port 37 nsew signal output
rlabel metal2 s 6458 200 6514 800 6 chanx_left_out[15]
port 38 nsew signal output
rlabel metal3 s 29200 21088 29800 21208 6 chanx_left_out[16]
port 39 nsew signal output
rlabel metal2 s 27710 200 27766 800 6 chanx_left_out[17]
port 40 nsew signal output
rlabel metal3 s 29200 10888 29800 11008 6 chanx_left_out[18]
port 41 nsew signal output
rlabel metal2 s 16118 29200 16174 29800 6 chanx_left_out[1]
port 42 nsew signal output
rlabel metal2 s 10322 29200 10378 29800 6 chanx_left_out[2]
port 43 nsew signal output
rlabel metal3 s 29200 8 29800 128 6 chanx_left_out[3]
port 44 nsew signal output
rlabel metal3 s 29200 22448 29800 22568 6 chanx_left_out[4]
port 45 nsew signal output
rlabel metal2 s 28998 29200 29054 29800 6 chanx_left_out[5]
port 46 nsew signal output
rlabel metal3 s 200 4768 800 4888 6 chanx_left_out[6]
port 47 nsew signal output
rlabel metal2 s 10322 200 10378 800 6 chanx_left_out[7]
port 48 nsew signal output
rlabel metal3 s 29200 4768 29800 4888 6 chanx_left_out[8]
port 49 nsew signal output
rlabel metal3 s 200 17008 800 17128 6 chanx_left_out[9]
port 50 nsew signal output
rlabel metal3 s 200 2048 800 2168 6 chany_bottom_in[0]
port 51 nsew signal input
rlabel metal3 s 200 23128 800 23248 6 chany_bottom_in[10]
port 52 nsew signal input
rlabel metal2 s 7746 29200 7802 29800 6 chany_bottom_in[11]
port 53 nsew signal input
rlabel metal2 s 21914 200 21970 800 6 chany_bottom_in[12]
port 54 nsew signal input
rlabel metal2 s 26422 29200 26478 29800 6 chany_bottom_in[13]
port 55 nsew signal input
rlabel metal2 s 18694 200 18750 800 6 chany_bottom_in[14]
port 56 nsew signal input
rlabel metal2 s 1950 200 2006 800 6 chany_bottom_in[15]
port 57 nsew signal input
rlabel metal3 s 200 14288 800 14408 6 chany_bottom_in[16]
port 58 nsew signal input
rlabel metal2 s 26422 200 26478 800 6 chany_bottom_in[17]
port 59 nsew signal input
rlabel metal3 s 29200 12248 29800 12368 6 chany_bottom_in[18]
port 60 nsew signal input
rlabel metal3 s 29200 7488 29800 7608 6 chany_bottom_in[1]
port 61 nsew signal input
rlabel metal2 s 20626 200 20682 800 6 chany_bottom_in[2]
port 62 nsew signal input
rlabel metal3 s 200 25848 800 25968 6 chany_bottom_in[3]
port 63 nsew signal input
rlabel metal3 s 29200 1368 29800 1488 6 chany_bottom_in[4]
port 64 nsew signal input
rlabel metal2 s 3882 29200 3938 29800 6 chany_bottom_in[5]
port 65 nsew signal input
rlabel metal3 s 29200 9528 29800 9648 6 chany_bottom_in[6]
port 66 nsew signal input
rlabel metal3 s 200 12248 800 12368 6 chany_bottom_in[7]
port 67 nsew signal input
rlabel metal2 s 23202 200 23258 800 6 chany_bottom_in[8]
port 68 nsew signal input
rlabel metal3 s 29200 19728 29800 19848 6 chany_bottom_in[9]
port 69 nsew signal input
rlabel metal2 s 13542 200 13598 800 6 chany_bottom_out[0]
port 70 nsew signal output
rlabel metal3 s 200 18368 800 18488 6 chany_bottom_out[10]
port 71 nsew signal output
rlabel metal2 s 14830 200 14886 800 6 chany_bottom_out[11]
port 72 nsew signal output
rlabel metal2 s 18 200 74 800 6 chany_bottom_out[12]
port 73 nsew signal output
rlabel metal2 s 17406 200 17462 800 6 chany_bottom_out[13]
port 74 nsew signal output
rlabel metal3 s 200 6128 800 6248 6 chany_bottom_out[14]
port 75 nsew signal output
rlabel metal2 s 14830 29200 14886 29800 6 chany_bottom_out[15]
port 76 nsew signal output
rlabel metal3 s 200 9528 800 9648 6 chany_bottom_out[16]
port 77 nsew signal output
rlabel metal2 s 662 29200 718 29800 6 chany_bottom_out[17]
port 78 nsew signal output
rlabel metal2 s 4526 200 4582 800 6 chany_bottom_out[18]
port 79 nsew signal output
rlabel metal2 s 662 200 718 800 6 chany_bottom_out[1]
port 80 nsew signal output
rlabel metal2 s 27710 29200 27766 29800 6 chany_bottom_out[2]
port 81 nsew signal output
rlabel metal2 s 20626 29200 20682 29800 6 chany_bottom_out[3]
port 82 nsew signal output
rlabel metal2 s 12898 200 12954 800 6 chany_bottom_out[4]
port 83 nsew signal output
rlabel metal2 s 29642 29200 29698 29800 6 chany_bottom_out[5]
port 84 nsew signal output
rlabel metal3 s 29200 2048 29800 2168 6 chany_bottom_out[6]
port 85 nsew signal output
rlabel metal3 s 200 6808 800 6928 6 chany_bottom_out[7]
port 86 nsew signal output
rlabel metal3 s 29200 15648 29800 15768 6 chany_bottom_out[8]
port 87 nsew signal output
rlabel metal2 s 5814 200 5870 800 6 chany_bottom_out[9]
port 88 nsew signal output
rlabel metal2 s 9034 200 9090 800 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 89 nsew signal input
rlabel metal3 s 200 10888 800 11008 6 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 90 nsew signal input
rlabel metal3 s 29200 17008 29800 17128 6 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 91 nsew signal input
rlabel metal2 s 16118 200 16174 800 6 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 92 nsew signal input
rlabel metal2 s 23846 29200 23902 29800 6 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 93 nsew signal input
rlabel metal2 s 23202 29200 23258 29800 6 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 94 nsew signal input
rlabel metal2 s 1950 29200 2006 29800 6 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 95 nsew signal input
rlabel metal2 s 6458 29200 6514 29800 6 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 96 nsew signal input
rlabel metal2 s 19338 200 19394 800 6 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 97 nsew signal input
rlabel metal3 s 200 8168 800 8288 6 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 98 nsew signal input
rlabel metal3 s 200 27208 800 27328 6 pReset
port 99 nsew signal input
rlabel metal3 s 29200 13608 29800 13728 6 prog_clk
port 100 nsew signal input
rlabel metal4 s 4417 2128 4737 27792 6 vccd1
port 101 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 27792 6 vccd1
port 101 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 27792 6 vccd1
port 101 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 27792 6 vccd1
port 101 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 27792 6 vssd1
port 102 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 27792 6 vssd1
port 102 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 27792 6 vssd1
port 102 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 27792 6 vssd1
port 102 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2116052
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/sb_4__4_/runs/22_12_30_10_32/results/signoff/sb_4__4_.magic.gds
string GDS_START 126516
<< end >>

