* NGSPICE file created from sb_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

.subckt sb_1__1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
+ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9]
+ chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13]
+ chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[1] chany_top_in[2]
+ chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7]
+ chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11]
+ chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16]
+ chany_top_out[17] chany_top_out[18] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
+ pReset prog_clk right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
+ vccd1 vssd1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1270_ net13 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_1
X_0985_ _0160_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
X_1606_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out _0449_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1468_ mux_bottom_track_1.INVTX1_4_.out _0311_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1399_ mux_bottom_track_1.INVTX1_1_.out _0242_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_8
X_1537_ mux_left_track_9.INVTX1_9_.out _0380_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ mem_top_track_16.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
X_1253_ net30 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1322_ net55 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1184_ clknet_4_4_0_prog_clk mem_left_track_9.DFFR_4_.Q _0106_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0968_ _0159_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__inv_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0899_ net28 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0822_ net67 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_9_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0684_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__inv_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0753_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1305_ net63 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1167_ clknet_4_3_0_prog_clk mem_bottom_track_25.DFFR_5_.Q _0089_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1098_ clknet_4_5_0_prog_clk mem_top_track_16.DFFR_2_.Q _0020_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1021_ _0152_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__buf_4
X_0805_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_0.out sky130_fd_sc_hd__inv_2
X_0667_ mem_bottom_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__inv_2
X_0736_ mem_top_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__inv_2
X_0598_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XFILLER_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1219_ clknet_4_10_0_prog_clk mem_bottom_track_33.DFFR_3_.Q _0141_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1570_ mux_left_track_25.INVTX1_10_.out _0413_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_8
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0521_ mem_bottom_track_1.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__inv_2
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 mux_bottom_track_33.INVTX1_4_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1004_ _0162_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__inv_2
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0719_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__inv_2
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1622_ mux_bottom_track_33.INVTX1_3_.out _0465_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0504_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__inv_2
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1553_ mux_left_track_17.INVTX1_9_.out _0396_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ mux_bottom_track_9.INVTX1_4_.out _0327_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0984_ _0160_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__inv_2
X_1605_ mux_bottom_track_33.INVTX1_0_.out _0448_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1536_ net185 _0379_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1467_ mux_bottom_track_1.INVTX1_8_.out _0310_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1398_ mux_left_track_1.INVTX1_9_.out _0241_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1252_ mux_left_track_33.out vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1321_ mux_top_track_8.out vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1183_ clknet_4_9_0_prog_clk mem_left_track_9.DFFR_5_.Q _0105_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0967_ _0159_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__inv_2
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1519_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out _0362_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_0898_ net34 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0752_ mem_top_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__inv_2
X_0821_ net25 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0683_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
X_1304_ net73 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1166_ clknet_4_1_0_prog_clk mem_bottom_track_25.DFFR_6_.Q _0088_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1097_ clknet_4_12_0_prog_clk mem_top_track_16.DFFR_3_.Q _0019_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1020_ _0163_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__inv_2
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0735_ mem_top_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__inv_2
X_0804_ net94 vssd1 vssd1 vccd1 vccd1 mux_top_track_24.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_1504__183 vssd1 vssd1 vccd1 vccd1 net183 _1504__183/LO sky130_fd_sc_hd__conb_1
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0666_ mem_bottom_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__inv_2
X_0597_ mem_left_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__inv_2
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1218_ clknet_4_10_0_prog_clk mem_bottom_track_33.DFFR_4_.Q _0140_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1149_ clknet_4_15_0_prog_clk mem_bottom_track_1.DFFR_0_.D _0071_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0520_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _0162_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__inv_2
XFILLER_30_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0718_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__inv_2
X_0649_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__inv_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1621_ net191 _0464_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1552_ net186 _0395_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0503_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1483_ mux_bottom_track_9.INVTX1_8_.out _0326_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0983_ _0160_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__inv_2
X_1604_ mux_left_track_33.INVTX1_5_.out _0447_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1535_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out _0378_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1397_ mux_left_track_1.INVTX1_8_.out _0240_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1466_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out _0309_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1320_ net57 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1251_ net32 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
X_1182_ clknet_4_12_0_prog_clk mem_left_track_9.DFFR_6_.Q _0104_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0966_ _0153_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__buf_4
X_0897_ net18 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1449_ mux_bottom_track_25.INVTX1_2_.out _0292_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1518_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out _0361_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0820_ net40 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0751_ mem_top_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__inv_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1303_ net74 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
X_0682_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__inv_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1096_ clknet_4_8_0_prog_clk mem_top_track_16.DFFR_4_.Q _0018_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1165_ clknet_4_10_0_prog_clk mem_bottom_track_17.DFFR_0_.D _0087_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_0949_ _0157_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
XFILLER_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0665_ mem_bottom_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__inv_2
X_0803_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_24.out sky130_fd_sc_hd__inv_2
X_0734_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__inv_2
X_0596_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__inv_2
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1148_ clknet_4_15_0_prog_clk mem_bottom_track_1.DFFR_0_.Q _0070_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1079_ clknet_4_10_0_prog_clk mem_top_track_0.DFFR_5_.Q _0001_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1217_ clknet_4_1_0_prog_clk mem_right_track_24.DFFR_7_.Q _0139_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_7 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1002_ _0162_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__inv_2
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0717_ mem_right_track_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
X_0648_ mem_bottom_track_9.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__inv_2
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0579_ mem_left_track_9.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__inv_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1620_ mux_left_track_33.INVTX1_7_.out _0463_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_1
X_0502_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__inv_2
X_1551_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out _0394_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1482_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out _0325_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0982_ _0160_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1603_ mux_bottom_track_33.INVTX1_6_.out _0446_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1465_ mux_bottom_track_1.INVTX1_3_.out _0308_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1534_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out _0377_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1396_ mux_left_track_1.INVTX1_7_.out _0239_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1250_ net33 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_2
X_1181_ clknet_4_10_0_prog_clk mem_bottom_track_33.DFFR_5_.Q _0103_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0896_ net20 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0965_ _0158_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__inv_2
X_1517_ mux_bottom_track_25.INVTX1_0_.out _0360_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1448_ mux_left_track_25.INVTX1_2_.out _0291_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1379_ mux_bottom_track_25.INVTX1_10_.out _0222_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0681_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__inv_2
X_0750_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__inv_2
X_1392__176 vssd1 vssd1 vccd1 vccd1 net176 _1392__176/LO sky130_fd_sc_hd__conb_1
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1302_ mux_bottom_track_9.out vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1095_ clknet_4_2_0_prog_clk mem_top_track_16.DFFR_5_.Q _0017_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1164_ clknet_4_3_0_prog_clk mem_bottom_track_17.DFFR_0_.Q _0086_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_0948_ _0157_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
X_0879_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_17.out sky130_fd_sc_hd__inv_2
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0802_ net93 vssd1 vssd1 vccd1 vccd1 mux_top_track_16.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0664_ mem_bottom_track_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__inv_2
X_0733_ mem_top_track_24.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
XFILLER_37_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0595_ mem_left_track_1.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__inv_2
X_1216_ clknet_4_1_0_prog_clk mem_right_track_32.DFFR_0_.Q _0138_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1078_ clknet_4_10_0_prog_clk mem_top_track_0.DFFR_6_.Q _0000_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1147_ clknet_4_14_0_prog_clk mem_bottom_track_1.DFFR_1_.Q _0069_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_8 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1001_ _0162_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__inv_2
X_0578_ mem_left_track_17.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__inv_2
X_0647_ mem_bottom_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
X_0716_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__inv_2
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0501_ mem_left_track_33.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__inv_2
X_1550_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out _0393_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1481_ mux_bottom_track_9.INVTX1_3_.out _0324_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0981_ _0160_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__inv_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1602_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out _0445_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1395_ mux_bottom_track_1.INVTX1_11_.out _0238_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1533_ mux_bottom_track_1.INVTX1_0_.out _0376_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1464_ mux_bottom_track_1.INVTX1_2_.out _0307_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ clknet_4_3_0_prog_clk mem_left_track_1.DFFR_0_.Q _0102_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0964_ _0158_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__inv_2
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1516_ mux_bottom_track_25.INVTX1_4_.out _0359_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0895_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_33.out sky130_fd_sc_hd__inv_2
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1378_ mux_bottom_track_9.INVTX1_10_.out _0221_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1447_ mux_bottom_track_25.INVTX1_1_.out _0290_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0680_ mem_right_track_24.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__inv_2
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1301_ net76 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1094_ clknet_4_10_0_prog_clk mem_top_track_16.DFFR_6_.Q _0016_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1163_ clknet_4_7_0_prog_clk mem_bottom_track_17.DFFR_1_.Q _0085_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_0947_ _0157_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
XFILLER_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0878_ net85 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0801_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_16.out sky130_fd_sc_hd__inv_2
X_0732_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
X_0663_ mem_bottom_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__inv_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0594_ mem_left_track_1.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__inv_2
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1215_ clknet_4_3_0_prog_clk mem_right_track_32.DFFR_1_.Q _0137_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_1146_ clknet_4_12_0_prog_clk mem_bottom_track_1.DFFR_2_.Q _0068_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1077_ _0153_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__inv_2
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1000_ _0162_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__inv_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0715_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__inv_2
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0646_ mem_bottom_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
X_0577_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__inv_2
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1129_ clknet_4_14_0_prog_clk mem_right_track_16.DFFR_3_.Q _0051_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0500_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
X_1480_ mux_bottom_track_9.INVTX1_2_.out _0323_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0629_ mem_bottom_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__inv_2
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0980_ _0160_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__inv_2
XFILLER_16_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1601_ mux_left_track_17.INVTX1_2_.out _0444_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1532_ mux_bottom_track_1.INVTX1_3_.out _0375_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_8_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1394_ mux_bottom_track_1.INVTX1_9_.out _0237_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1463_ mux_bottom_track_1.INVTX1_1_.out _0306_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0894_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_32.out sky130_fd_sc_hd__inv_2
X_0963_ _0158_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__inv_2
X_1515_ mux_bottom_track_25.INVTX1_8_.out _0358_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1377_ mux_bottom_track_25.INVTX1_9_.out _0220_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1446_ mux_left_track_25.INVTX1_8_.out _0289_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1300_ net77 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1162_ clknet_4_4_0_prog_clk mem_bottom_track_17.DFFR_2_.Q _0084_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1093_ clknet_4_2_0_prog_clk mem_top_track_0.DFFR_7_.Q _0015_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1440__179 vssd1 vssd1 vccd1 vccd1 net179 _1440__179/LO sky130_fd_sc_hd__conb_1
X_0946_ _0157_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0877_ net72 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_1429_ mux_left_track_17.INVTX1_8_.out _0272_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0731_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
X_0800_ net92 vssd1 vssd1 vccd1 vccd1 mux_top_track_8.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0662_ mem_bottom_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__inv_2
X_0593_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1214_ clknet_4_2_0_prog_clk mem_right_track_32.DFFR_2_.Q _0136_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
X_1145_ clknet_4_13_0_prog_clk mem_bottom_track_1.DFFR_3_.Q _0067_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1076_ _0153_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__inv_2
X_0929_ _0155_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__inv_2
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0714_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__inv_2
X_0645_ mem_bottom_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__inv_2
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0576_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
X_1059_ _0167_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__inv_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1128_ clknet_4_9_0_prog_clk mem_right_track_16.DFFR_4_.Q _0050_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0628_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0559_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__inv_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1462_ mux_bottom_track_1.INVTX1_7_.out _0305_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1600_ mux_bottom_track_33.INVTX1_1_.out _0443_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1531_ mux_left_track_1.INVTX1_8_.out _0374_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1393_ mux_bottom_track_1.INVTX1_8_.out _0236_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0893_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_32.out sky130_fd_sc_hd__inv_2
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0962_ _0158_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__inv_2
X_1445_ mux_left_track_25.INVTX1_7_.out _0288_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1514_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out _0357_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1376_ net175 _0219_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1472__181 vssd1 vssd1 vccd1 vccd1 net181 _1472__181/LO sky130_fd_sc_hd__conb_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1092_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_0_.Q _0014_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1161_ clknet_4_6_0_prog_clk mem_bottom_track_17.DFFR_3_.Q _0083_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0876_ net54 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0945_ _0157_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1428_ mux_left_track_17.INVTX1_7_.out _0271_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1359_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out _0202_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0661_ mem_bottom_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__inv_2
X_0730_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0592_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__inv_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1213_ clknet_4_9_0_prog_clk mem_right_track_32.DFFR_3_.Q _0135_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_32.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1075_ _0168_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__inv_2
X_1144_ clknet_4_15_0_prog_clk mem_bottom_track_1.DFFR_4_.Q _0066_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0859_ net38 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0928_ _0155_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__inv_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0713_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__inv_2
X_0644_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
X_0575_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__inv_2
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1058_ _0167_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__inv_2
X_1127_ clknet_4_11_0_prog_clk mem_right_track_16.DFFR_5_.Q _0049_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0558_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__inv_2
X_0627_ mem_bottom_track_17.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__inv_2
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1392_ net176 _0235_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1461_ mux_bottom_track_1.INVTX1_6_.out _0304_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1530_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out _0373_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0961_ _0158_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__inv_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0892_ net83 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_11_.out sky130_fd_sc_hd__inv_2
X_1444_ mux_left_track_9.INVTX1_8_.out _0287_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1513_ mux_bottom_track_25.INVTX1_3_.out _0356_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1375_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out _0218_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1091_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_1_.Q _0013_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_2
X_1160_ clknet_4_12_0_prog_clk mem_bottom_track_17.DFFR_4_.Q _0082_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0944_ _0153_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__buf_4
XFILLER_20_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0875_ net56 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1427_ mux_bottom_track_17.INVTX1_11_.out _0270_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1358_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out _0201_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1289_ net70 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0660_ mem_bottom_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__inv_2
X_0591_ mem_left_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1212_ clknet_4_12_0_prog_clk mem_right_track_32.DFFR_4_.Q _0134_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1074_ _0168_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__inv_2
X_1143_ clknet_4_13_0_prog_clk mem_bottom_track_1.DFFR_5_.Q _0065_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0927_ _0155_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__inv_2
X_0858_ net26 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0789_ mem_top_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__inv_2
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0574_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__inv_2
X_0643_ mem_bottom_track_9.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0712_ mem_right_track_8.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__inv_2
X_1126_ clknet_4_14_0_prog_clk mem_right_track_16.DFFR_6_.Q _0048_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1057_ _0167_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__inv_2
XFILLER_56_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0557_ mem_left_track_17.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
X_0626_ mem_bottom_track_17.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__inv_2
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1109_ clknet_4_10_0_prog_clk mem_top_track_16.DFFR_7_.Q _0031_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1391_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out _0234_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1460_ mux_bottom_track_1.INVTX1_5_.out _0303_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0609_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__inv_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ mux_bottom_track_33.INVTX1_3_.out _0432_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0960_ _0158_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
X_1512_ mux_bottom_track_25.INVTX1_2_.out _0355_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_0891_ net65 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_1443_ mux_bottom_track_25.INVTX1_10_.out _0286_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1374_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out _0217_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1090_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_2_.Q _0012_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1520__184 vssd1 vssd1 vccd1 vccd1 net184 _1520__184/LO sky130_fd_sc_hd__conb_1
X_0943_ _0156_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
X_0874_ net61 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_9_.out sky130_fd_sc_hd__inv_2
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1288_ net71 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
X_1426_ mux_bottom_track_17.INVTX1_9_.out _0269_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1357_ mux_top_track_8.INVTX1_0_.out _0200_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0590_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__inv_2
X_1211_ clknet_4_5_0_prog_clk mem_top_track_24.DFFR_7_.Q _0133_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1142_ clknet_4_13_0_prog_clk mem_bottom_track_1.DFFR_6_.Q _0064_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_1.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1073_ _0168_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__inv_2
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0857_ net33 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0926_ _0155_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__inv_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0788_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
X_1409_ mux_bottom_track_9.INVTX1_8_.out _0252_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0711_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__inv_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0573_ mem_left_track_9.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__inv_2
X_0642_ mem_bottom_track_17.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__inv_2
XFILLER_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1125_ clknet_4_7_0_prog_clk mem_right_track_0.DFFR_7_.Q _0047_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1056_ _0167_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__inv_2
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0909_ net86 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__buf_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0625_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__inv_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0556_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1108_ clknet_4_14_0_prog_clk mem_top_track_24.DFFR_0_.Q _0030_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1039_ _0165_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__inv_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1390_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out _0233_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1588_ mux_bottom_track_33.INVTX1_2_.out _0431_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0608_ mem_bottom_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__inv_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ mem_top_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__inv_2
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0890_ net57 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1511_ mux_bottom_track_25.INVTX1_1_.out _0354_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1442_ mux_bottom_track_25.INVTX1_9_.out _0285_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1373_ mux_top_track_16.INVTX1_0_.out _0216_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0873_ net49 vssd1 vssd1 vccd1 vccd1 mux_left_track_9.INVTX1_10_.out sky130_fd_sc_hd__inv_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0942_ _0156_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
X_1425_ mux_bottom_track_17.INVTX1_8_.out _0268_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1287_ mux_right_track_0.out vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1356_ mux_bottom_track_9.INVTX1_6_.out _0199_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1072_ _0168_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1141_ clknet_4_14_0_prog_clk mem_right_track_16.DFFR_7_.Q _0063_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1210_ clknet_4_5_0_prog_clk mem_top_track_32.DFFR_0_.Q _0132_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0787_ mem_top_track_0.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__inv_2
X_0925_ _0155_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__inv_2
X_0856_ net2 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1408_ net177 _0251_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1339_ mux_bottom_track_1.INVTX1_8_.out _0182_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0710_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__inv_2
X_0641_ mem_bottom_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__inv_2
X_0572_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1055_ _0167_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__inv_2
X_1124_ clknet_4_1_0_prog_clk mem_right_track_8.DFFR_0_.Q _0046_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0908_ net50 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0839_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_17.out sky130_fd_sc_hd__inv_2
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ mem_bottom_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__inv_2
XFILLER_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0555_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__inv_2
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1038_ _0165_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__inv_2
X_1107_ clknet_4_13_0_prog_clk mem_top_track_24.DFFR_1_.Q _0029_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0607_ mem_bottom_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0538_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__inv_2
X_1587_ mux_bottom_track_33.INVTX1_6_.out _0430_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1441_ mux_bottom_track_25.INVTX1_8_.out _0284_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1510_ mux_bottom_track_25.INVTX1_7_.out _0353_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1372_ mux_bottom_track_17.INVTX1_6_.out _0215_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0941_ _0156_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0872_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_9.out sky130_fd_sc_hd__inv_2
X_1424_ net178 _0267_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_2
X_1355_ mux_bottom_track_9.INVTX1_8_.out _0198_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1286_ net6 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1071_ _0168_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__inv_2
XFILLER_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1140_ clknet_4_13_0_prog_clk mem_right_track_24.DFFR_0_.Q _0062_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0924_ _0155_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__inv_2
X_0855_ net19 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0786_ mem_top_track_0.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__inv_2
X_1338_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out _0181_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1407_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out _0250_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_61_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1269_ net14 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0571_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__inv_2
X_0640_ mem_bottom_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__inv_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1054_ _0152_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__buf_4
X_1123_ clknet_4_2_0_prog_clk mem_right_track_8.DFFR_1_.Q _0045_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_0907_ net79 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0769_ mem_top_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__inv_2
X_0838_ net11 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0623_ mem_bottom_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__inv_2
X_0554_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__inv_2
XFILLER_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1106_ clknet_4_7_0_prog_clk mem_top_track_24.DFFR_2_.Q _0028_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1037_ _0165_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__inv_2
Xinput90 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ vssd1 vssd1 vccd1
+ vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ mux_left_track_33.INVTX1_6_.out _0429_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0606_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__inv_2
X_0537_ mem_top_track_32.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__inv_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1440_ net179 _0283_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1371_ mux_bottom_track_17.INVTX1_8_.out _0214_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ mux_left_track_25.INVTX1_9_.out _0412_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0940_ _0156_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0871_ net84 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_11_.out sky130_fd_sc_hd__inv_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1285_ net16 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_1
X_1423_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out _0266_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1354_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out _0197_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_51_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1488__182 vssd1 vssd1 vccd1 vccd1 net182 _1488__182/LO sky130_fd_sc_hd__conb_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1070_ _0168_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0854_ net7 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_9_.out sky130_fd_sc_hd__inv_2
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0923_ _0155_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
X_0785_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
X_1268_ mux_left_track_1.out vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
X_1337_ mux_bottom_track_17.INVTX1_4_.out _0180_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1406_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out _0249_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_61_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1199_ clknet_4_1_0_prog_clk mem_left_track_25.DFFR_5_.Q _0121_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0570_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__inv_2
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1122_ clknet_4_2_0_prog_clk mem_right_track_8.DFFR_2_.Q _0044_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1053_ _0166_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__inv_2
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0906_ net58 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0837_ net73 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0699_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__inv_2
X_0768_ mem_top_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__inv_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0622_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__inv_2
X_0553_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1105_ clknet_4_6_0_prog_clk mem_top_track_24.DFFR_3_.Q _0027_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1036_ _0165_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__inv_2
Xinput91 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ vssd1 vssd1 vccd1
+ vccd1 net91 sky130_fd_sc_hd__clkbuf_1
Xinput80 chany_top_in[8] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ net188 _0428_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__inv_2
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0605_ mem_bottom_track_25.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
X_1019_ _0163_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__inv_2
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1370_ mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out _0213_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_4_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1499_ mux_bottom_track_17.INVTX1_8_.out _0342_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_0519_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
X_1568_ net187 _0411_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0870_ net75 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1422_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out _0265_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
X_1284_ net17 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_1
X_1353_ mux_bottom_track_9.INVTX1_5_.out _0196_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0999_ _0152_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__buf_4
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0853_ net14 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_10_.out sky130_fd_sc_hd__inv_2
X_0922_ _0153_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__buf_4
X_1405_ mux_bottom_track_1.INVTX1_0_.out _0248_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_8
X_0784_ mem_top_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
Xinput1 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_ vssd1 vssd1 vccd1
+ vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_1336_ mux_bottom_track_1.INVTX1_4_.out _0179_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1267_ net25 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1198_ clknet_4_1_0_prog_clk mem_left_track_25.DFFR_6_.Q _0120_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0_prog_clk prog_clk vssd1 vssd1 vccd1 vccd1 clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1052_ _0166_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__inv_2
X_1121_ clknet_4_0_0_prog_clk mem_right_track_8.DFFR_3_.Q _0043_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0905_ net47 vssd1 vssd1 vccd1 vccd1 mux_left_track_33.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0767_ mem_top_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__inv_2
X_0836_ net80 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0698_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__inv_2
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ net58 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0621_ mem_bottom_track_17.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__inv_2
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0552_ mem_left_track_25.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__inv_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1035_ _0165_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__inv_2
X_1104_ clknet_4_7_0_prog_clk mem_top_track_24.DFFR_4_.Q _0026_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput81 chany_top_in[9] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_2
X_0819_ net29 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_5_.out sky130_fd_sc_hd__inv_2
Xinput70 chany_top_in[16] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput92 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ vssd1 vssd1 vccd1
+ vccd1 net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1584_ mux_bottom_track_33.INVTX1_7_.out _0427_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0604_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__inv_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0535_ mem_top_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1018_ _0163_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__inv_2
XFILLER_1_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0518_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
X_1567_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out _0410_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1498_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out _0341_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1421_ mux_bottom_track_9.INVTX1_0_.out _0264_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1352_ mux_bottom_track_9.INVTX1_4_.out _0195_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1283_ mux_right_track_8.out vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0998_ _0161_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__inv_2
X_1619_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out _0462_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_1536__185 vssd1 vssd1 vccd1 vccd1 net185 _1536__185/LO sky130_fd_sc_hd__conb_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ _0154_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__inv_2
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0783_ mem_top_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_0852_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1
+ vccd1 vccd1 mux_bottom_track_25.out sky130_fd_sc_hd__clkinv_2
X_1404_ mux_right_track_0.INVTX1_4_.out _0247_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1335_ mux_bottom_track_1.INVTX1_3_.out _0178_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1266_ net35 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_ vssd1 vssd1 vccd1
+ vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_1197_ clknet_4_14_0_prog_clk mem_left_track_17.DFFR_0_.D _0119_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1328__172 vssd1 vssd1 vccd1 vccd1 net172 _1328__172/LO sky130_fd_sc_hd__conb_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1120_ clknet_4_0_0_prog_clk mem_right_track_8.DFFR_4_.Q _0042_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1051_ _0166_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__inv_2
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0904_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_33.out sky130_fd_sc_hd__inv_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0697_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__inv_2
X_0766_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__inv_2
X_0835_ net68 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1318_ net59 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0620_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__inv_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0551_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1034_ _0165_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__inv_2
X_1103_ clknet_4_4_0_prog_clk mem_top_track_24.DFFR_5_.Q _0025_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput60 chany_bottom_in[7] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xinput93 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ vssd1 vssd1 vccd1
+ vccd1 net93 sky130_fd_sc_hd__clkbuf_1
Xinput82 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ vssd1 vssd1 vccd1
+ vccd1 net82 sky130_fd_sc_hd__clkbuf_1
X_0818_ net31 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0749_ mem_top_track_16.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__inv_2
Xinput71 chany_top_in[17] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0534_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__inv_2
X_1583_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out _0426_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0603_ mem_left_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
XFILLER_7_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1017_ _0163_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__inv_2
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1497_ mux_bottom_track_17.INVTX1_3_.out _0340_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1566_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out _0409_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_0517_ mem_right_track_32.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__inv_2
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1420_ mux_right_track_8.INVTX1_4_.out _0263_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1351_ mux_bottom_track_9.INVTX1_3_.out _0194_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1282_ net19 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1618_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out _0461_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_0997_ _0161_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__inv_2
X_1549_ mux_bottom_track_9.INVTX1_0_.out _0392_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0920_ _0154_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__inv_2
X_0851_ net13 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_11_.out sky130_fd_sc_hd__inv_2
X_0782_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
X_1403_ mux_left_track_33.INVTX1_7_.out _0246_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1265_ net36 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
X_1334_ mux_left_track_1.INVTX1_9_.out _0177_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
Xinput3 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_ vssd1 vssd1 vccd1
+ vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1196_ clknet_4_14_0_prog_clk mem_left_track_17.DFFR_0_.Q _0118_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1050_ _0166_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__inv_2
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0903_ net9 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0834_ net35 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0696_ mem_right_track_16.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
X_0765_ mem_top_track_8.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__inv_2
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1317_ mux_top_track_16.out vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ clknet_4_6_0_prog_clk mem_left_track_1.DFFR_1_.Q _0101_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 chany_top_out[8] sky130_fd_sc_hd__buf_2
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0550_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__inv_2
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1102_ clknet_4_4_0_prog_clk mem_top_track_24.DFFR_6_.Q _0024_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_24.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1033_ _0165_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__inv_2
Xinput50 chany_bottom_in[15] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
X_0817_ net3 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_7_.out sky130_fd_sc_hd__inv_2
Xinput61 chany_bottom_in[8] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 chany_top_in[18] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
X_0679_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__inv_2
X_0748_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
Xinput94 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_ vssd1 vssd1 vccd1
+ vccd1 net94 sky130_fd_sc_hd__clkbuf_1
Xinput83 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ vssd1 vssd1 vccd1
+ vccd1 net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out _0425_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0602_ mem_left_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__inv_2
X_0533_ mem_right_track_0.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__inv_2
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1016_ _0163_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__inv_2
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1565_ mux_bottom_track_17.INVTX1_0_.out _0408_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1496_ mux_bottom_track_17.INVTX1_2_.out _0339_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0516_ mem_bottom_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1281_ net20 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_2
X_1350_ mux_left_track_9.INVTX1_10_.out _0193_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0996_ _0161_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__inv_2
X_1617_ mux_bottom_track_33.INVTX1_0_.out _0460_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1479_ mux_bottom_track_9.INVTX1_1_.out _0322_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1548_ mux_bottom_track_9.INVTX1_3_.out _0391_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0850_ net74 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1402_ mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out _0245_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_0781_ mem_top_track_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
X_1264_ mux_left_track_9.out vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1333_ mux_left_track_1.INVTX1_8_.out _0176_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
Xinput4 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_ vssd1 vssd1 vccd1
+ vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1195_ clknet_4_15_0_prog_clk mem_left_track_17.DFFR_1_.Q _0117_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0979_ _0160_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__inv_2
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0902_ net77 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0833_ net42 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0695_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__inv_2
X_0764_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__inv_2
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1178_ clknet_4_2_0_prog_clk mem_left_track_1.DFFR_2_.Q _0100_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1316_ net61 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 chany_top_out[16] sky130_fd_sc_hd__buf_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 chany_top_out[9] sky130_fd_sc_hd__buf_2
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1032_ _0152_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__buf_4
X_1101_ clknet_4_0_0_prog_clk mem_top_track_16.DFFR_0_.D _0023_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput40 chanx_right_in[6] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dlymetal6s2s_1
X_0816_ net6 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0747_ mem_top_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__inv_2
Xinput73 chany_top_in[1] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_2
Xinput51 chany_bottom_in[16] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput62 chany_bottom_in[9] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ vssd1 vssd1 vccd1
+ vccd1 net84 sky130_fd_sc_hd__clkbuf_1
X_0678_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__inv_2
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1581_ mux_bottom_track_25.INVTX1_0_.out _0424_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_0601_ mem_left_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0532_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1015_ _0163_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__inv_2
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1564_ mux_bottom_track_17.INVTX1_3_.out _0407_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1495_ mux_bottom_track_17.INVTX1_1_.out _0338_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0515_ mem_bottom_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__inv_2
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1280_ net21 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0995_ _0161_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__inv_2
X_1547_ mux_left_track_9.INVTX1_8_.out _0390_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1616_ mux_bottom_track_33.INVTX1_3_.out _0459_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1478_ mux_bottom_track_9.INVTX1_7_.out _0321_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0780_ mem_top_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__inv_2
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1401_ mux_left_track_9.INVTX1_3_.out _0244_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_8
X_1263_ net38 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
X_1332_ mux_left_track_1.INVTX1_7_.out _0175_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1194_ clknet_4_11_0_prog_clk mem_left_track_17.DFFR_2_.Q _0116_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
Xinput5 ccff_head vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0978_ _0160_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__inv_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0901_ net66 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0763_ mem_top_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__inv_2
X_0832_ net27 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1315_ net62 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_1
X_0694_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1177_ clknet_4_9_0_prog_clk mem_left_track_1.DFFR_3_.Q _0099_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_10 mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 chany_top_out[17] sky130_fd_sc_hd__buf_2
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1100_ clknet_4_8_0_prog_clk mem_top_track_16.DFFR_0_.Q _0022_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1031_ _0164_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__inv_2
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput74 chany_top_in[2] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 chany_top_in[0] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dlymetal6s2s_1
X_0815_ net21 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0746_ mem_top_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__inv_2
Xinput85 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_ vssd1 vssd1 vccd1
+ vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xinput41 chanx_right_in[7] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
Xinput52 chany_bottom_in[17] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_2
Xinput30 chanx_right_in[14] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_2
X_0677_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__inv_2
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1229_ clknet_4_1_0_prog_clk mem_left_track_25.DFFR_7_.Q _0151_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0531_ mem_top_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__inv_2
X_1580_ mux_bottom_track_25.INVTX1_4_.out _0423_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0600_ mem_left_track_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__inv_2
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1014_ _0163_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__inv_2
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0729_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1563_ mux_left_track_17.INVTX1_8_.out _0406_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1494_ mux_bottom_track_17.INVTX1_7_.out _0337_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0514_ mem_bottom_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0994_ _0161_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__inv_2
X_1615_ mux_bottom_track_33.INVTX1_6_.out _0458_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1546_ mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out _0389_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1477_ mux_bottom_track_9.INVTX1_6_.out _0320_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1331_ mux_bottom_track_1.INVTX1_11_.out _0174_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1400_ mux_bottom_track_1.INVTX1_2_.out _0243_ vssd1 vssd1 vccd1 vccd1 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_8
Xinput6 chanx_left_in[0] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__dlymetal6s2s_1
X_1262_ net39 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
X_1193_ clknet_4_11_0_prog_clk mem_left_track_17.DFFR_3_.Q _0115_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0977_ _0153_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__buf_4
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1529_ mux_bottom_track_1.INVTX1_2_.out _0372_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0900_ net39 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0693_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__inv_2
X_0762_ mem_top_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
X_0831_ net30 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1314_ net45 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1176_ clknet_4_11_0_prog_clk mem_left_track_1.DFFR_4_.Q _0098_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_11 mem_top_track_0.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 chany_top_out[18] sky130_fd_sc_hd__buf_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[8] sky130_fd_sc_hd__buf_2
XFILLER_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1030_ _0164_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__inv_2
X_0814_ net22 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_10_.out sky130_fd_sc_hd__inv_2
Xinput31 chanx_right_in[15] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[5] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_2
Xinput64 chany_top_in[10] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 pReset vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
Xinput75 chany_top_in[3] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
X_0676_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__inv_2
Xinput53 chany_bottom_in[18] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
X_0745_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__inv_2
Xinput42 chanx_right_in[8] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1228_ clknet_4_3_0_prog_clk mem_left_track_33.DFFR_0_.Q _0150_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1159_ clknet_4_9_0_prog_clk mem_bottom_track_17.DFFR_5_.Q _0081_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0530_ mem_top_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__inv_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ _0163_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__inv_2
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0659_ mem_bottom_track_1.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__inv_2
X_0728_ mem_right_track_0.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__inv_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1493_ mux_bottom_track_17.INVTX1_6_.out _0336_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1562_ mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out _0405_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0513_ mem_bottom_track_33.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0993_ _0161_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__inv_2
X_1614_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out _0457_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1476_ mux_bottom_track_9.INVTX1_5_.out _0319_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1545_ mux_left_track_9.INVTX1_3_.out _0388_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1261_ net40 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_1
X_1330_ mux_bottom_track_1.INVTX1_9_.out _0173_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 chanx_left_in[10] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlymetal6s2s_1
X_1192_ clknet_4_11_0_prog_clk mem_left_track_17.DFFR_4_.Q _0114_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_0976_ _0159_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__inv_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1459_ mux_bottom_track_1.INVTX1_11_.out _0302_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1528_ mux_bottom_track_1.INVTX1_1_.out _0371_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0830_ net4 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0692_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__inv_2
X_0761_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
X_1313_ mux_top_track_24.out vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1175_ clknet_4_14_0_prog_clk mem_left_track_1.DFFR_5_.Q _0097_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_12 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0959_ _0158_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 chanx_right_out[6] sky130_fd_sc_hd__buf_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 chany_top_out[1] sky130_fd_sc_hd__buf_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[9] sky130_fd_sc_hd__buf_2
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 chanx_left_in[6] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
Xinput43 chanx_right_in[9] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dlymetal6s2s_1
X_0813_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_1.out sky130_fd_sc_hd__inv_2
Xinput54 chany_bottom_in[1] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_2
Xinput10 chanx_left_in[13] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 chanx_right_in[16] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_2
Xinput87 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ vssd1 vssd1 vccd1
+ vccd1 net87 sky130_fd_sc_hd__clkbuf_1
X_0744_ mem_top_track_24.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
X_0675_ mem_right_track_24.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__inv_2
Xinput76 chany_top_in[4] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput65 chany_top_in[11] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
X_1158_ clknet_4_11_0_prog_clk mem_bottom_track_17.DFFR_6_.Q _0080_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
X_1227_ clknet_4_4_0_prog_clk mem_left_track_33.DFFR_1_.Q _0149_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1089_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_3_.Q _0011_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ _0163_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__inv_2
X_0727_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__inv_2
XFILLER_57_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0658_ mem_bottom_track_1.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__inv_2
X_0589_ mem_left_track_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1492_ mux_bottom_track_17.INVTX1_5_.out _0335_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0512_ mem_bottom_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__inv_2
X_1561_ mux_bottom_track_17.INVTX1_2_.out _0404_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0992_ _0161_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__inv_2
X_1613_ mux_bottom_track_33.INVTX1_2_.out _0456_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1544_ mux_bottom_track_9.INVTX1_2_.out _0387_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1475_ mux_bottom_track_9.INVTX1_11_.out _0318_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[11] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_1191_ clknet_4_11_0_prog_clk mem_left_track_17.DFFR_5_.Q _0113_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1260_ mux_left_track_17.out vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0975_ _0159_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__inv_2
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1527_ mux_left_track_1.INVTX1_1_.out _0370_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1458_ mux_bottom_track_1.INVTX1_10_.out _0301_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1389_ mux_top_track_24.INVTX1_0_.out _0232_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ mem_top_track_16.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__inv_2
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0691_ mem_right_track_16.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__inv_2
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1312_ net47 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1174_ clknet_4_11_0_prog_clk mem_left_track_1.DFFR_6_.Q _0096_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_1.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0889_ net45 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0958_ _0158_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 chanx_right_out[7] sky130_fd_sc_hd__buf_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 chany_top_out[2] sky130_fd_sc_hd__buf_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput88 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ vssd1 vssd1 vccd1
+ vccd1 net88 sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_left_in[7] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 chanx_right_in[17] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_2
Xinput44 chany_bottom_in[0] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
X_0812_ net88 vssd1 vssd1 vccd1 vccd1 mux_right_track_24.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0743_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__inv_2
Xinput77 chany_top_in[5] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chanx_left_in[14] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput55 chany_bottom_in[2] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
Xinput66 chany_top_in[12] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_2
X_0674_ mem_right_track_24.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
X_1157_ clknet_4_9_0_prog_clk mem_bottom_track_1.DFFR_7_.Q _0079_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1226_ clknet_4_5_0_prog_clk mem_left_track_33.DFFR_2_.Q _0148_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1088_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_4_.Q _0010_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1011_ _0163_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__inv_2
XFILLER_19_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0726_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__inv_2
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0657_ mem_bottom_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__inv_2
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0588_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__inv_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1209_ clknet_4_4_0_prog_clk mem_top_track_32.DFFR_1_.Q _0131_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0511_ mem_bottom_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__inv_2
X_1560_ mux_left_track_17.INVTX1_2_.out _0403_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1491_ mux_bottom_track_17.INVTX1_11_.out _0334_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1552__186 vssd1 vssd1 vccd1 vccd1 net186 _1552__186/LO sky130_fd_sc_hd__conb_1
X_0709_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__inv_2
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1609__190 vssd1 vssd1 vccd1 vccd1 net190 _1609__190/LO sky130_fd_sc_hd__conb_1
X_0991_ _0161_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__inv_2
X_1612_ mux_bottom_track_33.INVTX1_1_.out _0455_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1474_ mux_bottom_track_9.INVTX1_10_.out _0317_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1543_ mux_bottom_track_9.INVTX1_1_.out _0386_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1344__173 vssd1 vssd1 vccd1 vccd1 net173 _1344__173/LO sky130_fd_sc_hd__conb_1
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1190_ clknet_4_10_0_prog_clk mem_left_track_17.DFFR_6_.Q _0112_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_17.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
Xinput9 chanx_left_in[12] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0974_ _0159_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__inv_2
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1457_ mux_bottom_track_1.INVTX1_9_.out _0300_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1526_ mux_left_track_1.INVTX1_7_.out _0369_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1388_ mux_bottom_track_33.INVTX1_4_.out _0231_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0690_ mem_right_track_16.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__inv_2
X_1311_ net48 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1173_ clknet_4_11_0_prog_clk mem_bottom_track_17.DFFR_7_.Q _0095_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 chanx_right_out[8] sky130_fd_sc_hd__buf_2
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_0888_ net46 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0957_ _0158_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 chany_top_out[10] sky130_fd_sc_hd__buf_2
X_1509_ mux_bottom_track_25.INVTX1_6_.out _0352_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 chany_top_out[3] sky130_fd_sc_hd__buf_2
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput56 chany_bottom_in[3] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
Xinput89 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_ vssd1 vssd1 vccd1
+ vccd1 net89 sky130_fd_sc_hd__clkbuf_1
X_0673_ mem_right_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__inv_2
X_0811_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_24.out sky130_fd_sc_hd__inv_2
X_0742_ mem_top_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
Xinput12 chanx_left_in[15] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 chanx_left_in[8] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_bottom_in[10] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput67 chany_top_in[13] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xinput34 chanx_right_in[18] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput78 chany_top_in[6] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1156_ clknet_4_3_0_prog_clk mem_bottom_track_9.DFFR_0_.Q _0078_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1087_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_5_.Q _0009_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_8.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1225_ clknet_4_5_0_prog_clk mem_left_track_33.DFFR_3_.Q _0147_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_33.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1010_ _0152_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__buf_4
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0725_ mem_right_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__inv_2
X_0656_ mem_bottom_track_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__inv_2
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1208_ clknet_4_4_0_prog_clk mem_top_track_32.DFFR_2_.Q _0130_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
X_0587_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
X_1585__188 vssd1 vssd1 vccd1 vccd1 net188 _1585__188/LO sky130_fd_sc_hd__conb_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1139_ clknet_4_12_0_prog_clk mem_right_track_24.DFFR_1_.Q _0061_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0510_ mem_bottom_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__inv_2
X_1490_ mux_bottom_track_17.INVTX1_10_.out _0333_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0708_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__inv_2
X_0639_ mem_bottom_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__inv_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1611_ mux_bottom_track_33.INVTX1_5_.out _0454_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0990_ _0161_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__inv_2
X_1473_ mux_bottom_track_9.INVTX1_9_.out _0316_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1542_ mux_left_track_9.INVTX1_7_.out _0385_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0973_ _0159_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__inv_2
X_1456_ net180 _0299_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1387_ mux_bottom_track_25.INVTX1_8_.out _0230_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1525_ mux_bottom_track_1.INVTX1_5_.out _0368_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1310_ net49 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1172_ clknet_4_15_0_prog_clk mem_bottom_track_25.DFFR_0_.Q _0094_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0956_ _0158_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 chany_top_out[11] sky130_fd_sc_hd__buf_2
X_0887_ net52 vssd1 vssd1 vccd1 vccd1 mux_left_track_25.INVTX1_10_.out sky130_fd_sc_hd__inv_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 chany_top_out[4] sky130_fd_sc_hd__buf_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 chanx_right_out[9] sky130_fd_sc_hd__buf_2
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1508_ mux_bottom_track_25.INVTX1_5_.out _0351_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1439_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out _0282_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput13 chanx_left_in[16] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dlymetal6s2s_1
X_0810_ net87 vssd1 vssd1 vccd1 vccd1 mux_right_track_16.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0741_ mem_top_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__inv_2
Xinput79 chany_top_in[7] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
Xinput57 chany_bottom_in[4] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_2
Xinput24 chanx_left_in[9] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 chanx_right_in[1] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput68 chany_top_in[14] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_2
Xinput46 chany_bottom_in[11] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0672_ mem_right_track_24.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__inv_2
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1224_ clknet_4_7_0_prog_clk mem_left_track_33.DFFR_4_.Q _0146_ vssd1 vssd1 vccd1
+ vccd1 net95 sky130_fd_sc_hd__dfrtp_2
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1155_ clknet_4_2_0_prog_clk mem_bottom_track_9.DFFR_1_.Q _0077_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_1086_ clknet_4_0_0_prog_clk mem_top_track_8.DFFR_6_.Q _0008_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_16.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0939_ _0156_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0724_ mem_right_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
X_0655_ mem_bottom_track_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__inv_2
X_0586_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__inv_2
X_1207_ clknet_4_4_0_prog_clk mem_top_track_32.DFFR_3_.Q _0129_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_32.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1069_ _0168_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__inv_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1138_ clknet_4_4_0_prog_clk mem_right_track_24.DFFR_2_.Q _0060_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0707_ mem_right_track_8.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__inv_2
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0569_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
X_0638_ mem_bottom_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__inv_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1610_ mux_bottom_track_33.INVTX1_4_.out _0453_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1472_ net181 _0315_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_2
X_1541_ mux_bottom_track_9.INVTX1_6_.out _0384_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0972_ _0159_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__inv_2
X_1524_ mux_bottom_track_1.INVTX1_4_.out _0367_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1455_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out _0298_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1386_ mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out _0229_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1171_ clknet_4_13_0_prog_clk mem_bottom_track_25.DFFR_1_.Q _0093_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0886_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_25.out sky130_fd_sc_hd__inv_2
X_0955_ _0153_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__buf_6
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 chany_top_out[5] sky130_fd_sc_hd__buf_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 chanx_right_out[17] sky130_fd_sc_hd__buf_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 chany_top_out[12] sky130_fd_sc_hd__buf_2
X_1507_ mux_bottom_track_25.INVTX1_11_.out _0350_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 chanx_left_out[14] sky130_fd_sc_hd__buf_2
X_1438_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out _0281_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1369_ mux_bottom_track_1.INVTX1_6_.out _0212_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 chanx_left_in[17] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
X_0740_ mem_top_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__inv_2
Xinput36 chanx_right_in[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_right_in[0] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput47 chany_bottom_in[12] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 chany_top_in[15] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_0671_ mem_right_track_24.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__inv_2
Xinput58 chany_bottom_in[5] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1154_ clknet_4_2_0_prog_clk mem_bottom_track_9.DFFR_2_.Q _0076_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1223_ clknet_4_1_0_prog_clk mem_bottom_track_25.DFFR_7_.Q _0145_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1085_ clknet_4_10_0_prog_clk net5 _0007_ vssd1 vssd1 vccd1 vccd1 mem_top_track_0.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_0869_ net44 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0938_ _0156_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0723_ mem_right_track_0.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__inv_2
X_0654_ mem_bottom_track_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__inv_2
X_0585_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1137_ clknet_4_1_0_prog_clk mem_right_track_24.DFFR_3_.Q _0059_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_1206_ clknet_4_5_0_prog_clk mem_top_track_32.DFFR_4_.Q _0128_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1068_ _0168_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__inv_2
XFILLER_25_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0706_ mem_right_track_16.DFFR_0_.D vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0499_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0568_ mem_left_track_17.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__inv_2
X_0637_ mem_bottom_track_9.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__inv_2
XFILLER_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1540_ mux_bottom_track_9.INVTX1_4_.out _0383_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1471_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out _0314_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0971_ _0159_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__inv_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1454_ mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out _0297_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1523_ mux_left_track_1.INVTX1_11_.out _0366_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1385_ mux_bottom_track_25.INVTX1_6_.out _0228_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1170_ clknet_4_5_0_prog_clk mem_bottom_track_25.DFFR_2_.Q _0092_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0885_ net82 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_11_.out sky130_fd_sc_hd__inv_2
X_0954_ _0157_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 chanx_left_out[15] sky130_fd_sc_hd__buf_2
X_1437_ mux_bottom_track_17.INVTX1_0_.out _0280_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1506_ mux_bottom_track_25.INVTX1_10_.out _0349_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 chany_top_out[13] sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 chany_top_out[6] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1368_ mux_bottom_track_17.INVTX1_5_.out _0211_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1299_ net78 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_1
XFILLER_62_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 chanx_right_in[3] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 chanx_left_in[18] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput26 chanx_right_in[10] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
X_0670_ mem_right_track_24.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__inv_2
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 chany_bottom_in[13] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 chany_bottom_in[6] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1222_ clknet_4_2_0_prog_clk mem_bottom_track_33.DFFR_0_.Q _0144_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1084_ clknet_4_10_0_prog_clk mem_top_track_0.DFFR_0_.Q _0006_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
X_1153_ clknet_4_8_0_prog_clk mem_bottom_track_9.DFFR_3_.Q _0075_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0868_ net59 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0937_ _0156_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
X_0799_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_8.out sky130_fd_sc_hd__clkinv_2
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0722_ mem_right_track_0.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__inv_2
X_0653_ mem_bottom_track_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__inv_2
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0584_ mem_left_track_9.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__inv_2
X_1205_ clknet_4_11_0_prog_clk mem_left_track_17.DFFR_7_.Q _0127_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1136_ clknet_4_1_0_prog_clk mem_right_track_24.DFFR_4_.Q _0058_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1067_ _0168_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__inv_2
XFILLER_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0636_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
X_0705_ mem_right_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__inv_2
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0498_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__inv_2
X_0567_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__inv_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1119_ clknet_4_0_0_prog_clk mem_right_track_8.DFFR_5_.Q _0041_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_8.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1470_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out _0313_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0619_ mem_bottom_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
X_1599_ mux_left_track_1.INVTX1_10_.out _0442_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0970_ _0159_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__inv_2
X_1453_ mux_bottom_track_25.INVTX1_0_.out _0296_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1522_ mux_left_track_1.INVTX1_10_.out _0365_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1384_ mux_bottom_track_25.INVTX1_5_.out _0227_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 chanx_left_out[16] sky130_fd_sc_hd__buf_2
X_0884_ net69 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0953_ _0157_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 chany_top_out[7] sky130_fd_sc_hd__buf_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[11] sky130_fd_sc_hd__buf_2
X_1436_ mux_right_track_16.INVTX1_4_.out _0279_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
X_1505_ mux_bottom_track_25.INVTX1_9_.out _0348_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1367_ mux_bottom_track_17.INVTX1_3_.out _0210_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 chany_top_out[14] sky130_fd_sc_hd__buf_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1298_ mux_bottom_track_17.out vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput38 chanx_right_in[4] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_2
Xinput49 chany_bottom_in[14] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput16 chanx_left_in[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 chanx_right_in[11] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1221_ clknet_4_9_0_prog_clk mem_bottom_track_33.DFFR_1_.Q _0143_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1083_ clknet_4_8_0_prog_clk mem_top_track_0.DFFR_1_.Q _0005_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_0.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
X_1152_ clknet_4_8_0_prog_clk mem_bottom_track_9.DFFR_4_.Q _0074_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0936_ _0156_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0867_ net48 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0798_ net91 vssd1 vssd1 vccd1 vccd1 mux_top_track_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_1419_ mux_left_track_9.INVTX1_10_.out _0262_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0721_ mem_right_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
X_0652_ mem_bottom_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__inv_2
X_0583_ mem_left_track_9.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__inv_2
XFILLER_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1204_ clknet_4_8_0_prog_clk mem_left_track_25.DFFR_0_.Q _0126_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1066_ _0168_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__inv_2
X_1135_ clknet_4_4_0_prog_clk mem_right_track_24.DFFR_5_.Q _0057_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_0919_ _0154_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__inv_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0566_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__inv_2
X_0635_ mem_bottom_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
X_0704_ mem_right_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
X_0497_ net95 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__inv_2
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1118_ clknet_4_0_0_prog_clk mem_right_track_8.DFFR_6_.Q _0040_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
X_1049_ _0166_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__inv_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1568__187 vssd1 vssd1 vccd1 vccd1 net187 _1568__187/LO sky130_fd_sc_hd__conb_1
XFILLER_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1598_ mux_left_track_33.INVTX1_6_.out _0441_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_0618_ mem_bottom_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__inv_2
X_0549_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__inv_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1452_ mux_right_track_24.INVTX1_4_.out _0295_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1383_ mux_bottom_track_25.INVTX1_4_.out _0226_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1521_ mux_left_track_1.INVTX1_9_.out _0364_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0952_ _0157_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XFILLER_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 chanx_right_out[2] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[5] sky130_fd_sc_hd__buf_2
X_1504_ net183 _0347_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 chany_top_out[15] sky130_fd_sc_hd__buf_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[12] sky130_fd_sc_hd__buf_2
X_0883_ net55 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_1435_ mux_left_track_17.INVTX1_10_.out _0278_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1366_ mux_left_track_17.INVTX1_10_.out _0209_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1297_ net80 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 chanx_left_in[2] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 chanx_right_in[12] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput39 chanx_right_in[5] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1151_ clknet_4_10_0_prog_clk mem_bottom_track_9.DFFR_5_.Q _0073_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_9.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
X_1220_ clknet_4_10_0_prog_clk mem_bottom_track_33.DFFR_2_.Q _0142_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_33.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1082_ clknet_4_8_0_prog_clk mem_top_track_0.DFFR_2_.Q _0004_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_0.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0935_ _0156_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
X_0866_ net53 vssd1 vssd1 vccd1 vccd1 mux_left_track_1.INVTX1_10_.out sky130_fd_sc_hd__inv_2
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0797_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_top_track_0.out sky130_fd_sc_hd__inv_2
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1418_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out _0261_ vssd1 vssd1
+ vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
X_1349_ mux_left_track_9.INVTX1_9_.out _0192_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0720_ mem_right_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__inv_2
X_0582_ mem_left_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__inv_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0651_ mem_bottom_track_9.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1203_ clknet_4_8_0_prog_clk mem_left_track_25.DFFR_1_.Q _0125_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1134_ clknet_4_6_0_prog_clk mem_right_track_24.DFFR_6_.Q _0056_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_24.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1065_ _0152_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__buf_4
X_0849_ net81 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0918_ _0154_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__inv_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0703_ mem_right_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__inv_2
X_0496_ mem_left_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__inv_2
X_0634_ mem_bottom_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
X_0565_ mem_left_track_17.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1117_ clknet_4_7_0_prog_clk mem_right_track_0.DFFR_0_.D _0039_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1048_ _0166_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__inv_2
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0617_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__inv_2
X_0548_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__inv_2
X_1597_ net189 _0440_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_53_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1520_ net184 _0363_ vssd1 vssd1 vccd1 vccd1 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1451_ mux_left_track_25.INVTX1_10_.out _0294_ vssd1 vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1382_ mux_left_track_25.INVTX1_10_.out _0225_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0882_ net60 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0951_ _0157_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 chanx_right_out[10] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1503_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out _0346_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 chanx_right_out[3] sky130_fd_sc_hd__buf_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 chanx_left_out[18] sky130_fd_sc_hd__buf_2
X_1296_ net81 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1365_ mux_left_track_17.INVTX1_9_.out _0208_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1434_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out _0277_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 chanx_left_in[3] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput29 chanx_right_in[13] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_1150_ clknet_4_10_0_prog_clk mem_bottom_track_9.DFFR_6_.Q _0072_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_17.DFFR_0_.D sky130_fd_sc_hd__dfrtp_1
X_1081_ clknet_4_8_0_prog_clk mem_top_track_0.DFFR_3_.Q _0003_ vssd1 vssd1 vccd1 vccd1
+ mem_top_track_0.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0865_ mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_left_track_1.out sky130_fd_sc_hd__inv_2
X_0934_ _0156_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0796_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__inv_2
X_1417_ mux_bottom_track_9.INVTX1_2_.out _0260_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1279_ mux_right_track_16.out vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_1
X_1348_ mux_left_track_9.INVTX1_7_.out _0191_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0650_ mem_bottom_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0581_ mem_left_track_9.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__inv_2
X_1064_ _0167_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__inv_2
X_1202_ clknet_4_8_0_prog_clk mem_left_track_25.DFFR_2_.Q _0124_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
X_1133_ clknet_4_6_0_prog_clk mem_right_track_16.DFFR_0_.D _0055_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0848_ net70 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0917_ _0154_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__inv_2
X_0779_ mem_top_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0702_ mem_right_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
X_0633_ mem_bottom_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__inv_2
X_0495_ mem_left_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
X_0564_ mem_left_track_17.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
X_1047_ _0166_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__inv_2
X_1116_ clknet_4_5_0_prog_clk mem_right_track_0.DFFR_0_.Q _0038_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1360__174 vssd1 vssd1 vccd1 vccd1 net174 _1360__174/LO sky130_fd_sc_hd__conb_1
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1596_ mux_bottom_track_33.INVTX1_7_.out _0439_ vssd1 vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_0616_ mem_bottom_track_25.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0547_ mem_left_track_25.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1450_ mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out _0293_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1381_ mux_left_track_25.INVTX1_8_.out _0224_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1408__177 vssd1 vssd1 vccd1 vccd1 net177 _1408__177/LO sky130_fd_sc_hd__conb_1
X_1579_ mux_left_track_25.INVTX1_8_.out _0422_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0881_ net62 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_9_.out sky130_fd_sc_hd__inv_2
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0950_ _0157_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 chanx_right_out[11] sky130_fd_sc_hd__buf_2
X_1433_ mux_bottom_track_17.INVTX1_2_.out _0276_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1502_ mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out _0345_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 chanx_right_out[4] sky130_fd_sc_hd__buf_2
X_1295_ net64 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_1
X_1364_ mux_left_track_17.INVTX1_7_.out _0207_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 chanx_left_in[4] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1080_ clknet_4_10_0_prog_clk mem_top_track_0.DFFR_4_.Q _0002_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_0.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0864_ net15 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_11_.out sky130_fd_sc_hd__inv_2
X_0795_ mem_top_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__inv_2
X_0933_ _0153_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__buf_4
X_1347_ mux_bottom_track_25.INVTX1_11_.out _0190_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1416_ mux_bottom_track_9.INVTX1_1_.out _0259_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1278_ net23 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0580_ mem_left_track_9.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__inv_2
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1201_ clknet_4_0_0_prog_clk mem_left_track_25.DFFR_3_.Q _0123_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_1063_ _0167_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__inv_2
X_1132_ clknet_4_13_0_prog_clk mem_right_track_16.DFFR_0_.Q _0054_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0916_ _0154_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
X_0847_ net36 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0778_ mem_top_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0632_ mem_bottom_track_17.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__inv_2
X_0701_ mem_right_track_8.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__inv_2
X_0563_ mem_left_track_17.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
X_0494_ mem_left_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1046_ _0166_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__inv_2
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1115_ clknet_4_6_0_prog_clk mem_right_track_0.DFFR_1_.Q _0037_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0615_ mem_bottom_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
X_0546_ mem_left_track_25.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__inv_2
X_1595_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out _0438_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1029_ _0164_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__inv_2
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1380_ mux_left_track_25.INVTX1_7_.out _0223_ vssd1 vssd1 vccd1 vccd1 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ mem_top_track_32.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__inv_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out _0421_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 chanx_left_out[2] sky130_fd_sc_hd__buf_2
X_0880_ net51 vssd1 vssd1 vccd1 vccd1 mux_left_track_17.INVTX1_10_.out sky130_fd_sc_hd__inv_2
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1432_ mux_bottom_track_17.INVTX1_1_.out _0275_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 chanx_right_out[12] sky130_fd_sc_hd__buf_2
X_1501_ mux_bottom_track_17.INVTX1_0_.out _0344_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1363_ mux_bottom_track_17.INVTX1_11_.out _0206_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 chanx_right_out[5] sky130_fd_sc_hd__buf_2
X_1294_ mux_bottom_track_25.out vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ _0155_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0863_ net76 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0794_ mem_top_track_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
X_1415_ mux_left_track_1.INVTX1_1_.out _0258_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1346_ mux_bottom_track_9.INVTX1_11_.out _0189_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1277_ net24 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1200_ clknet_4_0_0_prog_clk mem_left_track_25.DFFR_4_.Q _0122_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_25.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1062_ _0167_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__inv_2
X_1131_ clknet_4_5_0_prog_clk mem_right_track_16.DFFR_1_.Q _0053_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0915_ _0154_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0846_ net41 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0777_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__inv_2
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1329_ mux_bottom_track_33.INVTX1_5_.out _0172_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__inv_2
X_0631_ mem_bottom_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__inv_2
X_0562_ mem_left_track_17.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0493_ mem_left_track_33.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__inv_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1114_ clknet_4_1_0_prog_clk mem_right_track_0.DFFR_2_.Q _0036_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1045_ _0166_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__inv_2
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0829_ net16 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_8_.out sky130_fd_sc_hd__inv_2
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0614_ mem_bottom_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
X_0545_ mem_left_track_25.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__inv_2
X_1594_ mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out _0437_ vssd1
+ vssd1 vccd1 vccd1 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1028_ _0164_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__inv_2
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1577_ mux_bottom_track_25.INVTX1_2_.out _0420_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 chanx_left_out[3] sky130_fd_sc_hd__buf_2
X_1500_ mux_bottom_track_17.INVTX1_4_.out _0343_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1431_ mux_left_track_33.INVTX1_1_.out _0274_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1293_ net66 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
X_1362_ mux_bottom_track_17.INVTX1_10_.out _0205_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1629_ mux_bottom_track_33.INVTX1_0_.out _0472_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0862_ net64 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0931_ _0155_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0793_ mem_top_track_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
X_1276_ net7 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1345_ mux_bottom_track_9.INVTX1_9_.out _0188_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1414_ mux_left_track_25.INVTX1_9_.out _0257_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1130_ clknet_4_13_0_prog_clk mem_right_track_16.DFFR_2_.Q _0052_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_16.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1061_ _0167_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__inv_2
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0845_ net43 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_0914_ _0154_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__inv_2
X_0776_ mem_top_track_8.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
XFILLER_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1328_ net172 _0171_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1259_ net42 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0561_ mem_left_track_17.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
X_0630_ mem_bottom_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1044_ _0166_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__inv_2
X_1113_ clknet_4_1_0_prog_clk mem_right_track_0.DFFR_3_.Q _0035_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0759_ mem_top_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__inv_2
X_0828_ net23 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_9_.out sky130_fd_sc_hd__inv_2
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0613_ mem_bottom_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__inv_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ mux_bottom_track_25.INVTX1_3_.out _0436_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
X_0544_ mem_left_track_25.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1027_ _0164_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__inv_2
XFILLER_19_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1576_ mux_left_track_25.INVTX1_2_.out _0419_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_0527_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 chanx_left_out[4] sky130_fd_sc_hd__buf_2
X_1430_ mux_left_track_17.INVTX1_9_.out _0273_ vssd1 vssd1 vccd1 vccd1 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1361_ mux_bottom_track_17.INVTX1_9_.out _0204_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1292_ net67 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1559_ mux_bottom_track_17.INVTX1_1_.out _0402_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
X_1628_ mux_bottom_track_33.INVTX1_2_.out _0471_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0861_ net71 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_2_.out sky130_fd_sc_hd__inv_2
X_0930_ _0155_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__inv_2
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0792_ mem_top_track_0.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__inv_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1413_ mux_left_track_9.INVTX1_9_.out _0256_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1275_ mux_right_track_24.out vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1344_ net173 _0187_ vssd1 vssd1 vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1060_ _0167_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__inv_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0844_ net32 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_6_.out sky130_fd_sc_hd__inv_2
X_0775_ mem_top_track_8.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__inv_2
X_0913_ _0154_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__inv_2
X_1258_ net43 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
X_1189_ clknet_4_9_0_prog_clk mem_left_track_1.DFFR_7_.Q _0111_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
X_1327_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out _0170_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_17_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0560_ mem_left_track_17.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1043_ _0152_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__buf_6
X_1112_ clknet_4_7_0_prog_clk mem_right_track_0.DFFR_4_.Q _0034_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0827_ net8 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.INVTX1_10_.out sky130_fd_sc_hd__inv_2
X_0758_ mem_top_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
X_0689_ mem_right_track_16.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__inv_2
XFILLER_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0612_ mem_bottom_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__inv_2
X_1592_ mux_left_track_33.INVTX1_5_.out _0435_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0543_ mem_left_track_25.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1026_ _0164_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__inv_2
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0526_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
X_1575_ mux_bottom_track_25.INVTX1_1_.out _0418_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1009_ _0162_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1360_ net174 _0203_ vssd1 vssd1 vccd1 vccd1 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1291_ net68 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1627_ mux_left_track_33.INVTX1_6_.out _0470_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_1
X_1489_ mux_bottom_track_17.INVTX1_9_.out _0332_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
X_1558_ mux_left_track_17.INVTX1_7_.out _0401_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0509_ mem_bottom_track_33.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0860_ net37 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_25.INVTX1_3_.out sky130_fd_sc_hd__inv_2
X_0791_ mem_top_track_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__inv_2
X_1412_ mux_left_track_9.INVTX1_7_.out _0255_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1343_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out _0186_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
X_1274_ net9 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0989_ _0161_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__inv_2
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0912_ _0154_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
X_0843_ net1 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_7_.out sky130_fd_sc_hd__inv_2
X_0774_ mem_top_track_8.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
X_1326_ mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out _0169_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1188_ clknet_4_2_0_prog_clk mem_left_track_9.DFFR_0_.Q _0110_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_1_.Q sky130_fd_sc_hd__dfrtp_2
X_1257_ net26 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1042_ _0165_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__inv_2
X_1111_ clknet_4_7_0_prog_clk mem_right_track_0.DFFR_5_.Q _0033_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_6_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0688_ mem_right_track_16.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
X_0757_ mem_top_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__inv_2
X_0826_ mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_bottom_track_9.out sky130_fd_sc_hd__inv_2
X_1309_ mux_top_track_32.out vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ mux_bottom_track_1.INVTX1_10_.out _0434_ vssd1 vssd1 vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1376__175 vssd1 vssd1 vccd1 vccd1 net175 _1376__175/LO sky130_fd_sc_hd__conb_1
X_0542_ mem_left_track_25.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
X_0611_ mem_bottom_track_25.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__inv_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1025_ _0164_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__inv_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0809_ mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_16.out sky130_fd_sc_hd__inv_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_1 _0102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1574_ mux_left_track_25.INVTX1_7_.out _0417_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0525_ mem_right_track_32.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _0162_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__inv_2
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1290_ mux_bottom_track_33.out vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
X_1626_ mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out _0469_ vssd1 vssd1
+ vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0508_ mem_bottom_track_33.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
X_1557_ mux_bottom_track_17.INVTX1_6_.out _0400_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ net182 _0331_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0790_ mem_top_track_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__inv_2
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1273_ net10 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_1
X_1411_ mux_bottom_track_9.INVTX1_11_.out _0254_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1342_ mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out _0185_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0988_ _0153_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1609_ net190 _0452_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0842_ net17 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_8_.out sky130_fd_sc_hd__inv_2
X_0911_ _0153_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__buf_4
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0773_ mem_top_track_8.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__inv_2
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1256_ mux_left_track_25.out vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
X_1325_ mux_top_track_0.out vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_1
X_1187_ clknet_4_0_0_prog_clk mem_left_track_9.DFFR_1_.Q _0109_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1110_ clknet_4_13_0_prog_clk mem_right_track_0.DFFR_6_.Q _0032_ vssd1 vssd1 vccd1
+ vccd1 mem_right_track_0.DFFR_7_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ _0165_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__inv_2
X_0825_ net10 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_11_.out sky130_fd_sc_hd__inv_2
X_0756_ mem_top_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__inv_2
X_0687_ mem_right_track_16.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__inv_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1308_ net51 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out _0433_ vssd1 vssd1
+ vccd1 vccd1 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_0541_ mem_left_track_25.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__inv_2
X_0610_ mem_bottom_track_25.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1024_ _0164_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__inv_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0808_ net90 vssd1 vssd1 vccd1 vccd1 mux_right_track_8.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0739_ mem_top_track_24.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_2
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 mux_bottom_track_17.INVTX1_4_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1573_ mux_bottom_track_25.INVTX1_6_.out _0416_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_0524_ mem_right_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__inv_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1007_ _0162_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__inv_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1625_ mux_bottom_track_33.INVTX1_1_.out _0468_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1556_ mux_bottom_track_17.INVTX1_5_.out _0399_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0507_ mem_bottom_track_33.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
X_1487_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out _0330_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1410_ mux_bottom_track_9.INVTX1_9_.out _0253_ vssd1 vssd1 vccd1 vccd1 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1272_ net11 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1341_ mux_top_track_0.INVTX1_0_.out _0184_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0987_ _0160_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__inv_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1608_ mux_bottom_track_33.INVTX1_7_.out _0451_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1539_ mux_left_track_9.INVTX1_11_.out _0382_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0841_ net24 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_9_.out sky130_fd_sc_hd__inv_2
X_0910_ _0152_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_4
X_0772_ mem_top_track_8.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__inv_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1324_ net44 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
X_1255_ net28 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
X_1186_ clknet_4_2_0_prog_clk mem_left_track_9.DFFR_2_.Q _0108_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_3_.Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1040_ _0165_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__inv_2
X_0824_ net63 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_0_.out sky130_fd_sc_hd__inv_2
X_0755_ mem_top_track_16.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__inv_2
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0686_ mem_right_track_16.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__inv_2
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1307_ net52 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_1
X_1169_ clknet_4_4_0_prog_clk mem_bottom_track_25.DFFR_3_.Q _0091_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0540_ mem_top_track_32.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__inv_2
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1023_ _0164_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__inv_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1424__178 vssd1 vssd1 vccd1 vccd1 net178 _1424__178/LO sky130_fd_sc_hd__conb_1
X_0738_ mem_top_track_24.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__inv_2
X_0807_ mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out vssd1 vssd1 vccd1
+ vccd1 mux_right_track_8.out sky130_fd_sc_hd__clkinv_2
XFILLER_39_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0669_ mem_right_track_24.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__inv_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1572_ mux_bottom_track_25.INVTX1_5_.out _0415_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1597__189 vssd1 vssd1 vccd1 vccd1 net189 _1597__189/LO sky130_fd_sc_hd__conb_1
XANTENNA_3 mux_bottom_track_17.INVTX1_4_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0523_ mem_right_track_32.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1006_ _0162_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__inv_2
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1624_ mux_left_track_33.INVTX1_1_.out _0467_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_1
X_1555_ mux_left_track_17.INVTX1_11_.out _0398_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_0506_ mem_bottom_track_33.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__inv_2
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1486_ mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out _0329_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1340_ mux_bottom_track_1.INVTX1_5_.out _0183_ vssd1 vssd1 vccd1 vccd1 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
+ sky130_fd_sc_hd__ebufn_4
X_1271_ mux_right_track_32.out vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0986_ _0160_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__inv_2
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1469_ mux_bottom_track_1.INVTX1_0_.out _0312_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_2
X_1607_ mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out _0450_ vssd1
+ vssd1 vccd1 vccd1 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
+ sky130_fd_sc_hd__ebufn_4
X_1538_ mux_left_track_9.INVTX1_10_.out _0381_ vssd1 vssd1 vccd1 vccd1 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_4
XFILLER_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0840_ net12 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_17.INVTX1_10_.out sky130_fd_sc_hd__inv_2
X_0771_ mem_top_track_8.DFFR_6_.Q vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1323_ net54 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1254_ net29 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
X_1185_ clknet_4_0_0_prog_clk mem_left_track_9.DFFR_3_.Q _0107_ vssd1 vssd1 vccd1
+ vccd1 mem_left_track_9.DFFR_4_.Q sky130_fd_sc_hd__dfrtp_1
X_0969_ _0159_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__inv_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0823_ net78 vssd1 vssd1 vccd1 vccd1 mux_bottom_track_1.INVTX1_1_.out sky130_fd_sc_hd__inv_2
X_0685_ mem_right_track_16.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__inv_2
X_0754_ mem_top_track_16.DFFR_7_.Q vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__inv_2
X_1306_ mux_bottom_track_1.out vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1168_ clknet_4_6_0_prog_clk mem_bottom_track_25.DFFR_4_.Q _0090_ vssd1 vssd1 vccd1
+ vccd1 mem_bottom_track_25.DFFR_5_.Q sky130_fd_sc_hd__dfrtp_1
X_1099_ clknet_4_6_0_prog_clk mem_top_track_16.DFFR_1_.Q _0021_ vssd1 vssd1 vccd1
+ vccd1 mem_top_track_16.DFFR_2_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1456__180 vssd1 vssd1 vccd1 vccd1 net180 _1456__180/LO sky130_fd_sc_hd__conb_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1022_ _0164_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__inv_2
X_0806_ net89 vssd1 vssd1 vccd1 vccd1 mux_right_track_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_0737_ mem_top_track_24.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__inv_2
X_0668_ mem_bottom_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__inv_2
XFILLER_39_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0599_ mem_left_track_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0522_ mem_right_track_32.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 mux_bottom_track_33.INVTX1_4_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1571_ mux_left_track_25.INVTX1_11_.out _0414_ vssd1 vssd1 vccd1 vccd1 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_8
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1005_ _0162_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__inv_2
X_1621__191 vssd1 vssd1 vccd1 vccd1 net191 _1621__191/LO sky130_fd_sc_hd__conb_1
XFILLER_25_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1623_ mux_left_track_33.INVTX1_5_.out _0466_ vssd1 vssd1 vccd1 vccd1 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
X_1554_ mux_left_track_17.INVTX1_10_.out _0397_ vssd1 vssd1 vccd1 vccd1 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
+ sky130_fd_sc_hd__ebufn_2
X_1485_ mux_bottom_track_9.INVTX1_0_.out _0328_ vssd1 vssd1 vccd1 vccd1 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
+ sky130_fd_sc_hd__ebufn_4
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0505_ mem_bottom_track_33.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__inv_2
.ends

